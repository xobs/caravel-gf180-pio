VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_pio
  CLASS BLOCK ;
  FOREIGN wb_pio ;
  ORIGIN 0.000 0.000 ;
  SIZE 1300.000 BY 1400.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 1396.000 26.130 1400.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 1396.000 357.330 1400.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 1396.000 390.450 1400.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 1396.000 423.570 1400.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 1396.000 456.690 1400.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 1396.000 489.810 1400.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 1396.000 522.930 1400.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 1396.000 556.050 1400.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 1396.000 589.170 1400.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 1396.000 622.290 1400.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 1396.000 655.410 1400.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 1396.000 59.250 1400.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 1396.000 688.530 1400.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1396.000 721.650 1400.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 1396.000 754.770 1400.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 1396.000 787.890 1400.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 1396.000 821.010 1400.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.850 1396.000 854.130 1400.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 1396.000 887.250 1400.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.090 1396.000 920.370 1400.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1396.000 953.490 1400.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.330 1396.000 986.610 1400.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 1396.000 92.370 1400.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.450 1396.000 1019.730 1400.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 1396.000 1052.850 1400.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 1396.000 1085.970 1400.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 1396.000 1119.090 1400.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 1396.000 1152.210 1400.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 1396.000 1185.330 1400.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 1396.000 1218.450 1400.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.290 1396.000 1251.570 1400.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 1396.000 125.490 1400.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 1396.000 158.610 1400.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 1396.000 191.730 1400.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 1396.000 224.850 1400.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1396.000 257.970 1400.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 1396.000 291.090 1400.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 1396.000 324.210 1400.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 1396.000 37.170 1400.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 1396.000 368.370 1400.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 1396.000 401.490 1400.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 1396.000 434.610 1400.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 1396.000 467.730 1400.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 1396.000 500.850 1400.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 1396.000 533.970 1400.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 1396.000 567.090 1400.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 1396.000 600.210 1400.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 1396.000 633.330 1400.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 1396.000 666.450 1400.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 1396.000 70.290 1400.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 1396.000 699.570 1400.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 1396.000 732.690 1400.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 1396.000 765.810 1400.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 1396.000 798.930 1400.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 1396.000 832.050 1400.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 1396.000 865.170 1400.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 1396.000 898.290 1400.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 1396.000 931.410 1400.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 1396.000 964.530 1400.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.370 1396.000 997.650 1400.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 1396.000 103.410 1400.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 1396.000 1030.770 1400.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 1396.000 1063.890 1400.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.730 1396.000 1097.010 1400.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 1396.000 1130.130 1400.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.970 1396.000 1163.250 1400.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 1396.000 1196.370 1400.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.210 1396.000 1229.490 1400.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 1396.000 1262.610 1400.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 1396.000 136.530 1400.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 1396.000 169.650 1400.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 1396.000 202.770 1400.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 1396.000 235.890 1400.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 1396.000 269.010 1400.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 1396.000 302.130 1400.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 1396.000 335.250 1400.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 1396.000 48.210 1400.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 1396.000 379.410 1400.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 1396.000 412.530 1400.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 1396.000 445.650 1400.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 1396.000 478.770 1400.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 1396.000 511.890 1400.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 1396.000 545.010 1400.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 1396.000 578.130 1400.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 1396.000 611.250 1400.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 1396.000 644.370 1400.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 1396.000 677.490 1400.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 1396.000 81.330 1400.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 1396.000 710.610 1400.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 1396.000 743.730 1400.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 1396.000 776.850 1400.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 1396.000 809.970 1400.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 1396.000 843.090 1400.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 1396.000 876.210 1400.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.050 1396.000 909.330 1400.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.170 1396.000 942.450 1400.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 1396.000 975.570 1400.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 1396.000 1008.690 1400.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 1396.000 114.450 1400.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 1396.000 1041.810 1400.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.650 1396.000 1074.930 1400.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 1396.000 1108.050 1400.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 1396.000 1141.170 1400.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 1396.000 1174.290 1400.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.130 1396.000 1207.410 1400.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 1396.000 1240.530 1400.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.370 1396.000 1273.650 1400.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 1396.000 147.570 1400.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1396.000 180.690 1400.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 1396.000 213.810 1400.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 1396.000 246.930 1400.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 1396.000 280.050 1400.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 1396.000 313.170 1400.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 1396.000 346.290 1400.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 0.000 1213.390 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.410 0.000 1215.690 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.510 0.000 1024.790 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.410 0.000 1031.690 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.110 0.000 1052.390 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.010 0.000 1059.290 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 0.000 1066.190 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.810 0.000 1073.090 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.510 0.000 1093.790 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.410 0.000 1100.690 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.310 0.000 1107.590 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 0.000 1121.390 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.810 0.000 1142.090 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.710 0.000 1148.990 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 0.000 1155.890 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 0.000 1176.590 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.210 0.000 1183.490 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.110 0.000 1190.390 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.010 0.000 1197.290 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.910 0.000 1204.190 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.010 0.000 507.290 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 0.000 638.390 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 0.000 762.590 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 0.000 803.990 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 0.000 817.790 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 0.000 824.690 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 0.000 838.490 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 0.000 845.390 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 0.000 852.290 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.810 0.000 866.090 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 0.000 893.690 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 0.000 900.590 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.010 0.000 921.290 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 0.000 941.990 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.510 0.000 955.790 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.910 0.000 997.190 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.810 0.000 1004.090 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 0.000 1010.990 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 0.000 1020.190 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 0.000 1040.890 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 0.000 1047.790 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 0.000 1061.590 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 0.000 1068.490 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1088.910 0.000 1089.190 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 0.000 1123.690 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.310 0.000 1130.590 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.110 0.000 1144.390 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 0.000 1151.290 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 0.000 1158.190 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 0.000 1165.090 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.710 0.000 1171.990 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 0.000 1185.790 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 0.000 1192.690 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 0.000 1199.590 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 0.000 1206.490 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 0.000 757.990 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 0.000 778.690 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 0.000 799.390 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 0.000 813.190 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 0.000 826.990 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 0.000 833.890 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 0.000 861.490 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 0.000 868.390 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 0.000 882.190 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.310 0.000 923.590 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 0.000 937.390 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 0.000 958.090 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 0.000 978.790 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 0.000 985.690 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 0.000 999.490 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.110 0.000 1006.390 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 0.000 1022.490 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 0.000 1029.390 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.810 0.000 1050.090 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.710 0.000 1056.990 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 0.000 1084.590 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.010 0.000 1105.290 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 0.000 1112.190 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.810 0.000 1119.090 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.610 0.000 1132.890 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 0.000 1139.790 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.210 0.000 1160.490 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1167.110 0.000 1167.390 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.010 0.000 1174.290 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 0.000 1194.990 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 0.000 1201.890 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 0.000 767.190 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.810 0.000 774.090 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 0.000 836.190 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.110 0.000 891.390 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 0.000 912.090 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 0.000 918.990 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.310 0.000 946.590 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 0.000 967.290 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 0.000 974.190 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 0.000 1001.790 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 0.000 1015.590 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1387.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1387.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1387.440 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 1383.065 1294.630 1385.895 ;
        RECT 5.330 1377.625 1294.630 1380.455 ;
        RECT 5.330 1372.185 1294.630 1375.015 ;
        RECT 5.330 1366.745 1294.630 1369.575 ;
        RECT 5.330 1361.305 1294.630 1364.135 ;
        RECT 5.330 1355.865 1294.630 1358.695 ;
        RECT 5.330 1350.425 1294.630 1353.255 ;
        RECT 5.330 1344.985 1294.630 1347.815 ;
        RECT 5.330 1339.545 1294.630 1342.375 ;
        RECT 5.330 1334.105 1294.630 1336.935 ;
        RECT 5.330 1328.665 1294.630 1331.495 ;
        RECT 5.330 1323.225 1294.630 1326.055 ;
        RECT 5.330 1317.785 1294.630 1320.615 ;
        RECT 5.330 1312.345 1294.630 1315.175 ;
        RECT 5.330 1306.905 1294.630 1309.735 ;
        RECT 5.330 1301.465 1294.630 1304.295 ;
        RECT 5.330 1296.025 1294.630 1298.855 ;
        RECT 5.330 1290.585 1294.630 1293.415 ;
        RECT 5.330 1285.145 1294.630 1287.975 ;
        RECT 5.330 1279.705 1294.630 1282.535 ;
        RECT 5.330 1274.265 1294.630 1277.095 ;
        RECT 5.330 1268.825 1294.630 1271.655 ;
        RECT 5.330 1263.385 1294.630 1266.215 ;
        RECT 5.330 1257.945 1294.630 1260.775 ;
        RECT 5.330 1252.505 1294.630 1255.335 ;
        RECT 5.330 1247.065 1294.630 1249.895 ;
        RECT 5.330 1241.625 1294.630 1244.455 ;
        RECT 5.330 1236.185 1294.630 1239.015 ;
        RECT 5.330 1230.745 1294.630 1233.575 ;
        RECT 5.330 1225.305 1294.630 1228.135 ;
        RECT 5.330 1219.865 1294.630 1222.695 ;
        RECT 5.330 1214.425 1294.630 1217.255 ;
        RECT 5.330 1208.985 1294.630 1211.815 ;
        RECT 5.330 1203.545 1294.630 1206.375 ;
        RECT 5.330 1198.105 1294.630 1200.935 ;
        RECT 5.330 1192.665 1294.630 1195.495 ;
        RECT 5.330 1187.225 1294.630 1190.055 ;
        RECT 5.330 1181.785 1294.630 1184.615 ;
        RECT 5.330 1176.345 1294.630 1179.175 ;
        RECT 5.330 1170.905 1294.630 1173.735 ;
        RECT 5.330 1165.465 1294.630 1168.295 ;
        RECT 5.330 1160.025 1294.630 1162.855 ;
        RECT 5.330 1154.585 1294.630 1157.415 ;
        RECT 5.330 1149.145 1294.630 1151.975 ;
        RECT 5.330 1143.705 1294.630 1146.535 ;
        RECT 5.330 1138.265 1294.630 1141.095 ;
        RECT 5.330 1132.825 1294.630 1135.655 ;
        RECT 5.330 1127.385 1294.630 1130.215 ;
        RECT 5.330 1121.945 1294.630 1124.775 ;
        RECT 5.330 1116.505 1294.630 1119.335 ;
        RECT 5.330 1111.065 1294.630 1113.895 ;
        RECT 5.330 1105.625 1294.630 1108.455 ;
        RECT 5.330 1100.185 1294.630 1103.015 ;
        RECT 5.330 1094.745 1294.630 1097.575 ;
        RECT 5.330 1089.305 1294.630 1092.135 ;
        RECT 5.330 1083.865 1294.630 1086.695 ;
        RECT 5.330 1078.425 1294.630 1081.255 ;
        RECT 5.330 1072.985 1294.630 1075.815 ;
        RECT 5.330 1067.545 1294.630 1070.375 ;
        RECT 5.330 1062.105 1294.630 1064.935 ;
        RECT 5.330 1056.665 1294.630 1059.495 ;
        RECT 5.330 1051.225 1294.630 1054.055 ;
        RECT 5.330 1045.785 1294.630 1048.615 ;
        RECT 5.330 1040.345 1294.630 1043.175 ;
        RECT 5.330 1034.905 1294.630 1037.735 ;
        RECT 5.330 1029.465 1294.630 1032.295 ;
        RECT 5.330 1024.025 1294.630 1026.855 ;
        RECT 5.330 1018.585 1294.630 1021.415 ;
        RECT 5.330 1013.145 1294.630 1015.975 ;
        RECT 5.330 1007.705 1294.630 1010.535 ;
        RECT 5.330 1002.265 1294.630 1005.095 ;
        RECT 5.330 996.825 1294.630 999.655 ;
        RECT 5.330 991.385 1294.630 994.215 ;
        RECT 5.330 985.945 1294.630 988.775 ;
        RECT 5.330 980.505 1294.630 983.335 ;
        RECT 5.330 975.065 1294.630 977.895 ;
        RECT 5.330 969.625 1294.630 972.455 ;
        RECT 5.330 964.185 1294.630 967.015 ;
        RECT 5.330 958.745 1294.630 961.575 ;
        RECT 5.330 953.305 1294.630 956.135 ;
        RECT 5.330 947.865 1294.630 950.695 ;
        RECT 5.330 942.425 1294.630 945.255 ;
        RECT 5.330 936.985 1294.630 939.815 ;
        RECT 5.330 931.545 1294.630 934.375 ;
        RECT 5.330 926.105 1294.630 928.935 ;
        RECT 5.330 920.665 1294.630 923.495 ;
        RECT 5.330 915.225 1294.630 918.055 ;
        RECT 5.330 909.785 1294.630 912.615 ;
        RECT 5.330 904.345 1294.630 907.175 ;
        RECT 5.330 898.905 1294.630 901.735 ;
        RECT 5.330 893.465 1294.630 896.295 ;
        RECT 5.330 888.025 1294.630 890.855 ;
        RECT 5.330 882.585 1294.630 885.415 ;
        RECT 5.330 877.145 1294.630 879.975 ;
        RECT 5.330 871.705 1294.630 874.535 ;
        RECT 5.330 866.265 1294.630 869.095 ;
        RECT 5.330 860.825 1294.630 863.655 ;
        RECT 5.330 855.385 1294.630 858.215 ;
        RECT 5.330 849.945 1294.630 852.775 ;
        RECT 5.330 844.505 1294.630 847.335 ;
        RECT 5.330 839.065 1294.630 841.895 ;
        RECT 5.330 833.625 1294.630 836.455 ;
        RECT 5.330 828.185 1294.630 831.015 ;
        RECT 5.330 822.745 1294.630 825.575 ;
        RECT 5.330 817.305 1294.630 820.135 ;
        RECT 5.330 811.865 1294.630 814.695 ;
        RECT 5.330 806.425 1294.630 809.255 ;
        RECT 5.330 800.985 1294.630 803.815 ;
        RECT 5.330 795.545 1294.630 798.375 ;
        RECT 5.330 790.105 1294.630 792.935 ;
        RECT 5.330 784.665 1294.630 787.495 ;
        RECT 5.330 779.225 1294.630 782.055 ;
        RECT 5.330 773.785 1294.630 776.615 ;
        RECT 5.330 768.345 1294.630 771.175 ;
        RECT 5.330 762.905 1294.630 765.735 ;
        RECT 5.330 757.465 1294.630 760.295 ;
        RECT 5.330 752.025 1294.630 754.855 ;
        RECT 5.330 746.585 1294.630 749.415 ;
        RECT 5.330 741.145 1294.630 743.975 ;
        RECT 5.330 735.705 1294.630 738.535 ;
        RECT 5.330 730.265 1294.630 733.095 ;
        RECT 5.330 724.825 1294.630 727.655 ;
        RECT 5.330 719.385 1294.630 722.215 ;
        RECT 5.330 713.945 1294.630 716.775 ;
        RECT 5.330 708.505 1294.630 711.335 ;
        RECT 5.330 703.065 1294.630 705.895 ;
        RECT 5.330 697.625 1294.630 700.455 ;
        RECT 5.330 692.185 1294.630 695.015 ;
        RECT 5.330 686.745 1294.630 689.575 ;
        RECT 5.330 681.305 1294.630 684.135 ;
        RECT 5.330 675.865 1294.630 678.695 ;
        RECT 5.330 670.425 1294.630 673.255 ;
        RECT 5.330 664.985 1294.630 667.815 ;
        RECT 5.330 659.545 1294.630 662.375 ;
        RECT 5.330 654.105 1294.630 656.935 ;
        RECT 5.330 648.665 1294.630 651.495 ;
        RECT 5.330 643.225 1294.630 646.055 ;
        RECT 5.330 637.785 1294.630 640.615 ;
        RECT 5.330 632.345 1294.630 635.175 ;
        RECT 5.330 626.905 1294.630 629.735 ;
        RECT 5.330 621.465 1294.630 624.295 ;
        RECT 5.330 616.025 1294.630 618.855 ;
        RECT 5.330 610.585 1294.630 613.415 ;
        RECT 5.330 605.145 1294.630 607.975 ;
        RECT 5.330 599.705 1294.630 602.535 ;
        RECT 5.330 594.265 1294.630 597.095 ;
        RECT 5.330 588.825 1294.630 591.655 ;
        RECT 5.330 583.385 1294.630 586.215 ;
        RECT 5.330 577.945 1294.630 580.775 ;
        RECT 5.330 572.505 1294.630 575.335 ;
        RECT 5.330 567.065 1294.630 569.895 ;
        RECT 5.330 561.625 1294.630 564.455 ;
        RECT 5.330 556.185 1294.630 559.015 ;
        RECT 5.330 550.745 1294.630 553.575 ;
        RECT 5.330 545.305 1294.630 548.135 ;
        RECT 5.330 539.865 1294.630 542.695 ;
        RECT 5.330 534.425 1294.630 537.255 ;
        RECT 5.330 528.985 1294.630 531.815 ;
        RECT 5.330 523.545 1294.630 526.375 ;
        RECT 5.330 518.105 1294.630 520.935 ;
        RECT 5.330 512.665 1294.630 515.495 ;
        RECT 5.330 507.225 1294.630 510.055 ;
        RECT 5.330 501.785 1294.630 504.615 ;
        RECT 5.330 496.345 1294.630 499.175 ;
        RECT 5.330 490.905 1294.630 493.735 ;
        RECT 5.330 485.465 1294.630 488.295 ;
        RECT 5.330 480.025 1294.630 482.855 ;
        RECT 5.330 474.585 1294.630 477.415 ;
        RECT 5.330 469.145 1294.630 471.975 ;
        RECT 5.330 463.705 1294.630 466.535 ;
        RECT 5.330 458.265 1294.630 461.095 ;
        RECT 5.330 452.825 1294.630 455.655 ;
        RECT 5.330 447.385 1294.630 450.215 ;
        RECT 5.330 441.945 1294.630 444.775 ;
        RECT 5.330 436.505 1294.630 439.335 ;
        RECT 5.330 431.065 1294.630 433.895 ;
        RECT 5.330 425.625 1294.630 428.455 ;
        RECT 5.330 420.185 1294.630 423.015 ;
        RECT 5.330 414.745 1294.630 417.575 ;
        RECT 5.330 409.305 1294.630 412.135 ;
        RECT 5.330 403.865 1294.630 406.695 ;
        RECT 5.330 398.425 1294.630 401.255 ;
        RECT 5.330 392.985 1294.630 395.815 ;
        RECT 5.330 387.545 1294.630 390.375 ;
        RECT 5.330 382.105 1294.630 384.935 ;
        RECT 5.330 376.665 1294.630 379.495 ;
        RECT 5.330 371.225 1294.630 374.055 ;
        RECT 5.330 365.785 1294.630 368.615 ;
        RECT 5.330 360.345 1294.630 363.175 ;
        RECT 5.330 354.905 1294.630 357.735 ;
        RECT 5.330 349.465 1294.630 352.295 ;
        RECT 5.330 344.025 1294.630 346.855 ;
        RECT 5.330 338.585 1294.630 341.415 ;
        RECT 5.330 333.145 1294.630 335.975 ;
        RECT 5.330 327.705 1294.630 330.535 ;
        RECT 5.330 322.265 1294.630 325.095 ;
        RECT 5.330 316.825 1294.630 319.655 ;
        RECT 5.330 311.385 1294.630 314.215 ;
        RECT 5.330 305.945 1294.630 308.775 ;
        RECT 5.330 300.505 1294.630 303.335 ;
        RECT 5.330 295.065 1294.630 297.895 ;
        RECT 5.330 289.625 1294.630 292.455 ;
        RECT 5.330 284.185 1294.630 287.015 ;
        RECT 5.330 278.745 1294.630 281.575 ;
        RECT 5.330 273.305 1294.630 276.135 ;
        RECT 5.330 267.865 1294.630 270.695 ;
        RECT 5.330 262.425 1294.630 265.255 ;
        RECT 5.330 256.985 1294.630 259.815 ;
        RECT 5.330 251.545 1294.630 254.375 ;
        RECT 5.330 246.105 1294.630 248.935 ;
        RECT 5.330 240.665 1294.630 243.495 ;
        RECT 5.330 235.225 1294.630 238.055 ;
        RECT 5.330 229.785 1294.630 232.615 ;
        RECT 5.330 224.345 1294.630 227.175 ;
        RECT 5.330 218.905 1294.630 221.735 ;
        RECT 5.330 213.465 1294.630 216.295 ;
        RECT 5.330 208.025 1294.630 210.855 ;
        RECT 5.330 202.585 1294.630 205.415 ;
        RECT 5.330 197.145 1294.630 199.975 ;
        RECT 5.330 191.705 1294.630 194.535 ;
        RECT 5.330 186.265 1294.630 189.095 ;
        RECT 5.330 180.825 1294.630 183.655 ;
        RECT 5.330 175.385 1294.630 178.215 ;
        RECT 5.330 169.945 1294.630 172.775 ;
        RECT 5.330 164.505 1294.630 167.335 ;
        RECT 5.330 159.065 1294.630 161.895 ;
        RECT 5.330 153.625 1294.630 156.455 ;
        RECT 5.330 148.185 1294.630 151.015 ;
        RECT 5.330 142.745 1294.630 145.575 ;
        RECT 5.330 137.305 1294.630 140.135 ;
        RECT 5.330 131.865 1294.630 134.695 ;
        RECT 5.330 126.425 1294.630 129.255 ;
        RECT 5.330 120.985 1294.630 123.815 ;
        RECT 5.330 115.545 1294.630 118.375 ;
        RECT 5.330 110.105 1294.630 112.935 ;
        RECT 5.330 104.665 1294.630 107.495 ;
        RECT 5.330 99.225 1294.630 102.055 ;
        RECT 5.330 93.785 1294.630 96.615 ;
        RECT 5.330 88.345 1294.630 91.175 ;
        RECT 5.330 82.905 1294.630 85.735 ;
        RECT 5.330 77.465 1294.630 80.295 ;
        RECT 5.330 72.025 1294.630 74.855 ;
        RECT 5.330 66.585 1294.630 69.415 ;
        RECT 5.330 61.145 1294.630 63.975 ;
        RECT 5.330 55.705 1294.630 58.535 ;
        RECT 5.330 50.265 1294.630 53.095 ;
        RECT 5.330 44.825 1294.630 47.655 ;
        RECT 5.330 39.385 1294.630 42.215 ;
        RECT 5.330 33.945 1294.630 36.775 ;
        RECT 5.330 28.505 1294.630 31.335 ;
        RECT 5.330 23.065 1294.630 25.895 ;
        RECT 5.330 17.625 1294.630 20.455 ;
        RECT 5.330 12.185 1294.630 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1294.440 1387.285 ;
      LAYER met1 ;
        RECT 5.520 8.200 1294.440 1387.440 ;
      LAYER met2 ;
        RECT 8.380 1395.720 25.570 1396.450 ;
        RECT 26.410 1395.720 36.610 1396.450 ;
        RECT 37.450 1395.720 47.650 1396.450 ;
        RECT 48.490 1395.720 58.690 1396.450 ;
        RECT 59.530 1395.720 69.730 1396.450 ;
        RECT 70.570 1395.720 80.770 1396.450 ;
        RECT 81.610 1395.720 91.810 1396.450 ;
        RECT 92.650 1395.720 102.850 1396.450 ;
        RECT 103.690 1395.720 113.890 1396.450 ;
        RECT 114.730 1395.720 124.930 1396.450 ;
        RECT 125.770 1395.720 135.970 1396.450 ;
        RECT 136.810 1395.720 147.010 1396.450 ;
        RECT 147.850 1395.720 158.050 1396.450 ;
        RECT 158.890 1395.720 169.090 1396.450 ;
        RECT 169.930 1395.720 180.130 1396.450 ;
        RECT 180.970 1395.720 191.170 1396.450 ;
        RECT 192.010 1395.720 202.210 1396.450 ;
        RECT 203.050 1395.720 213.250 1396.450 ;
        RECT 214.090 1395.720 224.290 1396.450 ;
        RECT 225.130 1395.720 235.330 1396.450 ;
        RECT 236.170 1395.720 246.370 1396.450 ;
        RECT 247.210 1395.720 257.410 1396.450 ;
        RECT 258.250 1395.720 268.450 1396.450 ;
        RECT 269.290 1395.720 279.490 1396.450 ;
        RECT 280.330 1395.720 290.530 1396.450 ;
        RECT 291.370 1395.720 301.570 1396.450 ;
        RECT 302.410 1395.720 312.610 1396.450 ;
        RECT 313.450 1395.720 323.650 1396.450 ;
        RECT 324.490 1395.720 334.690 1396.450 ;
        RECT 335.530 1395.720 345.730 1396.450 ;
        RECT 346.570 1395.720 356.770 1396.450 ;
        RECT 357.610 1395.720 367.810 1396.450 ;
        RECT 368.650 1395.720 378.850 1396.450 ;
        RECT 379.690 1395.720 389.890 1396.450 ;
        RECT 390.730 1395.720 400.930 1396.450 ;
        RECT 401.770 1395.720 411.970 1396.450 ;
        RECT 412.810 1395.720 423.010 1396.450 ;
        RECT 423.850 1395.720 434.050 1396.450 ;
        RECT 434.890 1395.720 445.090 1396.450 ;
        RECT 445.930 1395.720 456.130 1396.450 ;
        RECT 456.970 1395.720 467.170 1396.450 ;
        RECT 468.010 1395.720 478.210 1396.450 ;
        RECT 479.050 1395.720 489.250 1396.450 ;
        RECT 490.090 1395.720 500.290 1396.450 ;
        RECT 501.130 1395.720 511.330 1396.450 ;
        RECT 512.170 1395.720 522.370 1396.450 ;
        RECT 523.210 1395.720 533.410 1396.450 ;
        RECT 534.250 1395.720 544.450 1396.450 ;
        RECT 545.290 1395.720 555.490 1396.450 ;
        RECT 556.330 1395.720 566.530 1396.450 ;
        RECT 567.370 1395.720 577.570 1396.450 ;
        RECT 578.410 1395.720 588.610 1396.450 ;
        RECT 589.450 1395.720 599.650 1396.450 ;
        RECT 600.490 1395.720 610.690 1396.450 ;
        RECT 611.530 1395.720 621.730 1396.450 ;
        RECT 622.570 1395.720 632.770 1396.450 ;
        RECT 633.610 1395.720 643.810 1396.450 ;
        RECT 644.650 1395.720 654.850 1396.450 ;
        RECT 655.690 1395.720 665.890 1396.450 ;
        RECT 666.730 1395.720 676.930 1396.450 ;
        RECT 677.770 1395.720 687.970 1396.450 ;
        RECT 688.810 1395.720 699.010 1396.450 ;
        RECT 699.850 1395.720 710.050 1396.450 ;
        RECT 710.890 1395.720 721.090 1396.450 ;
        RECT 721.930 1395.720 732.130 1396.450 ;
        RECT 732.970 1395.720 743.170 1396.450 ;
        RECT 744.010 1395.720 754.210 1396.450 ;
        RECT 755.050 1395.720 765.250 1396.450 ;
        RECT 766.090 1395.720 776.290 1396.450 ;
        RECT 777.130 1395.720 787.330 1396.450 ;
        RECT 788.170 1395.720 798.370 1396.450 ;
        RECT 799.210 1395.720 809.410 1396.450 ;
        RECT 810.250 1395.720 820.450 1396.450 ;
        RECT 821.290 1395.720 831.490 1396.450 ;
        RECT 832.330 1395.720 842.530 1396.450 ;
        RECT 843.370 1395.720 853.570 1396.450 ;
        RECT 854.410 1395.720 864.610 1396.450 ;
        RECT 865.450 1395.720 875.650 1396.450 ;
        RECT 876.490 1395.720 886.690 1396.450 ;
        RECT 887.530 1395.720 897.730 1396.450 ;
        RECT 898.570 1395.720 908.770 1396.450 ;
        RECT 909.610 1395.720 919.810 1396.450 ;
        RECT 920.650 1395.720 930.850 1396.450 ;
        RECT 931.690 1395.720 941.890 1396.450 ;
        RECT 942.730 1395.720 952.930 1396.450 ;
        RECT 953.770 1395.720 963.970 1396.450 ;
        RECT 964.810 1395.720 975.010 1396.450 ;
        RECT 975.850 1395.720 986.050 1396.450 ;
        RECT 986.890 1395.720 997.090 1396.450 ;
        RECT 997.930 1395.720 1008.130 1396.450 ;
        RECT 1008.970 1395.720 1019.170 1396.450 ;
        RECT 1020.010 1395.720 1030.210 1396.450 ;
        RECT 1031.050 1395.720 1041.250 1396.450 ;
        RECT 1042.090 1395.720 1052.290 1396.450 ;
        RECT 1053.130 1395.720 1063.330 1396.450 ;
        RECT 1064.170 1395.720 1074.370 1396.450 ;
        RECT 1075.210 1395.720 1085.410 1396.450 ;
        RECT 1086.250 1395.720 1096.450 1396.450 ;
        RECT 1097.290 1395.720 1107.490 1396.450 ;
        RECT 1108.330 1395.720 1118.530 1396.450 ;
        RECT 1119.370 1395.720 1129.570 1396.450 ;
        RECT 1130.410 1395.720 1140.610 1396.450 ;
        RECT 1141.450 1395.720 1151.650 1396.450 ;
        RECT 1152.490 1395.720 1162.690 1396.450 ;
        RECT 1163.530 1395.720 1173.730 1396.450 ;
        RECT 1174.570 1395.720 1184.770 1396.450 ;
        RECT 1185.610 1395.720 1195.810 1396.450 ;
        RECT 1196.650 1395.720 1206.850 1396.450 ;
        RECT 1207.690 1395.720 1217.890 1396.450 ;
        RECT 1218.730 1395.720 1228.930 1396.450 ;
        RECT 1229.770 1395.720 1239.970 1396.450 ;
        RECT 1240.810 1395.720 1251.010 1396.450 ;
        RECT 1251.850 1395.720 1262.050 1396.450 ;
        RECT 1262.890 1395.720 1273.090 1396.450 ;
        RECT 8.380 4.280 1273.640 1395.720 ;
        RECT 8.380 3.670 83.530 4.280 ;
        RECT 84.370 3.670 85.830 4.280 ;
        RECT 86.670 3.670 88.130 4.280 ;
        RECT 88.970 3.670 90.430 4.280 ;
        RECT 91.270 3.670 92.730 4.280 ;
        RECT 93.570 3.670 95.030 4.280 ;
        RECT 95.870 3.670 97.330 4.280 ;
        RECT 98.170 3.670 99.630 4.280 ;
        RECT 100.470 3.670 101.930 4.280 ;
        RECT 102.770 3.670 104.230 4.280 ;
        RECT 105.070 3.670 106.530 4.280 ;
        RECT 107.370 3.670 108.830 4.280 ;
        RECT 109.670 3.670 111.130 4.280 ;
        RECT 111.970 3.670 113.430 4.280 ;
        RECT 114.270 3.670 115.730 4.280 ;
        RECT 116.570 3.670 118.030 4.280 ;
        RECT 118.870 3.670 120.330 4.280 ;
        RECT 121.170 3.670 122.630 4.280 ;
        RECT 123.470 3.670 124.930 4.280 ;
        RECT 125.770 3.670 127.230 4.280 ;
        RECT 128.070 3.670 129.530 4.280 ;
        RECT 130.370 3.670 131.830 4.280 ;
        RECT 132.670 3.670 134.130 4.280 ;
        RECT 134.970 3.670 136.430 4.280 ;
        RECT 137.270 3.670 138.730 4.280 ;
        RECT 139.570 3.670 141.030 4.280 ;
        RECT 141.870 3.670 143.330 4.280 ;
        RECT 144.170 3.670 145.630 4.280 ;
        RECT 146.470 3.670 147.930 4.280 ;
        RECT 148.770 3.670 150.230 4.280 ;
        RECT 151.070 3.670 152.530 4.280 ;
        RECT 153.370 3.670 154.830 4.280 ;
        RECT 155.670 3.670 157.130 4.280 ;
        RECT 157.970 3.670 159.430 4.280 ;
        RECT 160.270 3.670 161.730 4.280 ;
        RECT 162.570 3.670 164.030 4.280 ;
        RECT 164.870 3.670 166.330 4.280 ;
        RECT 167.170 3.670 168.630 4.280 ;
        RECT 169.470 3.670 170.930 4.280 ;
        RECT 171.770 3.670 173.230 4.280 ;
        RECT 174.070 3.670 175.530 4.280 ;
        RECT 176.370 3.670 177.830 4.280 ;
        RECT 178.670 3.670 180.130 4.280 ;
        RECT 180.970 3.670 182.430 4.280 ;
        RECT 183.270 3.670 184.730 4.280 ;
        RECT 185.570 3.670 187.030 4.280 ;
        RECT 187.870 3.670 189.330 4.280 ;
        RECT 190.170 3.670 191.630 4.280 ;
        RECT 192.470 3.670 193.930 4.280 ;
        RECT 194.770 3.670 196.230 4.280 ;
        RECT 197.070 3.670 198.530 4.280 ;
        RECT 199.370 3.670 200.830 4.280 ;
        RECT 201.670 3.670 203.130 4.280 ;
        RECT 203.970 3.670 205.430 4.280 ;
        RECT 206.270 3.670 207.730 4.280 ;
        RECT 208.570 3.670 210.030 4.280 ;
        RECT 210.870 3.670 212.330 4.280 ;
        RECT 213.170 3.670 214.630 4.280 ;
        RECT 215.470 3.670 216.930 4.280 ;
        RECT 217.770 3.670 219.230 4.280 ;
        RECT 220.070 3.670 221.530 4.280 ;
        RECT 222.370 3.670 223.830 4.280 ;
        RECT 224.670 3.670 226.130 4.280 ;
        RECT 226.970 3.670 228.430 4.280 ;
        RECT 229.270 3.670 230.730 4.280 ;
        RECT 231.570 3.670 233.030 4.280 ;
        RECT 233.870 3.670 235.330 4.280 ;
        RECT 236.170 3.670 237.630 4.280 ;
        RECT 238.470 3.670 239.930 4.280 ;
        RECT 240.770 3.670 242.230 4.280 ;
        RECT 243.070 3.670 244.530 4.280 ;
        RECT 245.370 3.670 246.830 4.280 ;
        RECT 247.670 3.670 249.130 4.280 ;
        RECT 249.970 3.670 251.430 4.280 ;
        RECT 252.270 3.670 253.730 4.280 ;
        RECT 254.570 3.670 256.030 4.280 ;
        RECT 256.870 3.670 258.330 4.280 ;
        RECT 259.170 3.670 260.630 4.280 ;
        RECT 261.470 3.670 262.930 4.280 ;
        RECT 263.770 3.670 265.230 4.280 ;
        RECT 266.070 3.670 267.530 4.280 ;
        RECT 268.370 3.670 269.830 4.280 ;
        RECT 270.670 3.670 272.130 4.280 ;
        RECT 272.970 3.670 274.430 4.280 ;
        RECT 275.270 3.670 276.730 4.280 ;
        RECT 277.570 3.670 279.030 4.280 ;
        RECT 279.870 3.670 281.330 4.280 ;
        RECT 282.170 3.670 283.630 4.280 ;
        RECT 284.470 3.670 285.930 4.280 ;
        RECT 286.770 3.670 288.230 4.280 ;
        RECT 289.070 3.670 290.530 4.280 ;
        RECT 291.370 3.670 292.830 4.280 ;
        RECT 293.670 3.670 295.130 4.280 ;
        RECT 295.970 3.670 297.430 4.280 ;
        RECT 298.270 3.670 299.730 4.280 ;
        RECT 300.570 3.670 302.030 4.280 ;
        RECT 302.870 3.670 304.330 4.280 ;
        RECT 305.170 3.670 306.630 4.280 ;
        RECT 307.470 3.670 308.930 4.280 ;
        RECT 309.770 3.670 311.230 4.280 ;
        RECT 312.070 3.670 313.530 4.280 ;
        RECT 314.370 3.670 315.830 4.280 ;
        RECT 316.670 3.670 318.130 4.280 ;
        RECT 318.970 3.670 320.430 4.280 ;
        RECT 321.270 3.670 322.730 4.280 ;
        RECT 323.570 3.670 325.030 4.280 ;
        RECT 325.870 3.670 327.330 4.280 ;
        RECT 328.170 3.670 329.630 4.280 ;
        RECT 330.470 3.670 331.930 4.280 ;
        RECT 332.770 3.670 334.230 4.280 ;
        RECT 335.070 3.670 336.530 4.280 ;
        RECT 337.370 3.670 338.830 4.280 ;
        RECT 339.670 3.670 341.130 4.280 ;
        RECT 341.970 3.670 343.430 4.280 ;
        RECT 344.270 3.670 345.730 4.280 ;
        RECT 346.570 3.670 348.030 4.280 ;
        RECT 348.870 3.670 350.330 4.280 ;
        RECT 351.170 3.670 352.630 4.280 ;
        RECT 353.470 3.670 354.930 4.280 ;
        RECT 355.770 3.670 357.230 4.280 ;
        RECT 358.070 3.670 359.530 4.280 ;
        RECT 360.370 3.670 361.830 4.280 ;
        RECT 362.670 3.670 364.130 4.280 ;
        RECT 364.970 3.670 366.430 4.280 ;
        RECT 367.270 3.670 368.730 4.280 ;
        RECT 369.570 3.670 371.030 4.280 ;
        RECT 371.870 3.670 373.330 4.280 ;
        RECT 374.170 3.670 375.630 4.280 ;
        RECT 376.470 3.670 377.930 4.280 ;
        RECT 378.770 3.670 380.230 4.280 ;
        RECT 381.070 3.670 382.530 4.280 ;
        RECT 383.370 3.670 384.830 4.280 ;
        RECT 385.670 3.670 387.130 4.280 ;
        RECT 387.970 3.670 389.430 4.280 ;
        RECT 390.270 3.670 391.730 4.280 ;
        RECT 392.570 3.670 394.030 4.280 ;
        RECT 394.870 3.670 396.330 4.280 ;
        RECT 397.170 3.670 398.630 4.280 ;
        RECT 399.470 3.670 400.930 4.280 ;
        RECT 401.770 3.670 403.230 4.280 ;
        RECT 404.070 3.670 405.530 4.280 ;
        RECT 406.370 3.670 407.830 4.280 ;
        RECT 408.670 3.670 410.130 4.280 ;
        RECT 410.970 3.670 412.430 4.280 ;
        RECT 413.270 3.670 414.730 4.280 ;
        RECT 415.570 3.670 417.030 4.280 ;
        RECT 417.870 3.670 419.330 4.280 ;
        RECT 420.170 3.670 421.630 4.280 ;
        RECT 422.470 3.670 423.930 4.280 ;
        RECT 424.770 3.670 426.230 4.280 ;
        RECT 427.070 3.670 428.530 4.280 ;
        RECT 429.370 3.670 430.830 4.280 ;
        RECT 431.670 3.670 433.130 4.280 ;
        RECT 433.970 3.670 435.430 4.280 ;
        RECT 436.270 3.670 437.730 4.280 ;
        RECT 438.570 3.670 440.030 4.280 ;
        RECT 440.870 3.670 442.330 4.280 ;
        RECT 443.170 3.670 444.630 4.280 ;
        RECT 445.470 3.670 446.930 4.280 ;
        RECT 447.770 3.670 449.230 4.280 ;
        RECT 450.070 3.670 451.530 4.280 ;
        RECT 452.370 3.670 453.830 4.280 ;
        RECT 454.670 3.670 456.130 4.280 ;
        RECT 456.970 3.670 458.430 4.280 ;
        RECT 459.270 3.670 460.730 4.280 ;
        RECT 461.570 3.670 463.030 4.280 ;
        RECT 463.870 3.670 465.330 4.280 ;
        RECT 466.170 3.670 467.630 4.280 ;
        RECT 468.470 3.670 469.930 4.280 ;
        RECT 470.770 3.670 472.230 4.280 ;
        RECT 473.070 3.670 474.530 4.280 ;
        RECT 475.370 3.670 476.830 4.280 ;
        RECT 477.670 3.670 479.130 4.280 ;
        RECT 479.970 3.670 481.430 4.280 ;
        RECT 482.270 3.670 483.730 4.280 ;
        RECT 484.570 3.670 486.030 4.280 ;
        RECT 486.870 3.670 488.330 4.280 ;
        RECT 489.170 3.670 490.630 4.280 ;
        RECT 491.470 3.670 492.930 4.280 ;
        RECT 493.770 3.670 495.230 4.280 ;
        RECT 496.070 3.670 497.530 4.280 ;
        RECT 498.370 3.670 499.830 4.280 ;
        RECT 500.670 3.670 502.130 4.280 ;
        RECT 502.970 3.670 504.430 4.280 ;
        RECT 505.270 3.670 506.730 4.280 ;
        RECT 507.570 3.670 509.030 4.280 ;
        RECT 509.870 3.670 511.330 4.280 ;
        RECT 512.170 3.670 513.630 4.280 ;
        RECT 514.470 3.670 515.930 4.280 ;
        RECT 516.770 3.670 518.230 4.280 ;
        RECT 519.070 3.670 520.530 4.280 ;
        RECT 521.370 3.670 522.830 4.280 ;
        RECT 523.670 3.670 525.130 4.280 ;
        RECT 525.970 3.670 527.430 4.280 ;
        RECT 528.270 3.670 529.730 4.280 ;
        RECT 530.570 3.670 532.030 4.280 ;
        RECT 532.870 3.670 534.330 4.280 ;
        RECT 535.170 3.670 536.630 4.280 ;
        RECT 537.470 3.670 538.930 4.280 ;
        RECT 539.770 3.670 541.230 4.280 ;
        RECT 542.070 3.670 543.530 4.280 ;
        RECT 544.370 3.670 545.830 4.280 ;
        RECT 546.670 3.670 548.130 4.280 ;
        RECT 548.970 3.670 550.430 4.280 ;
        RECT 551.270 3.670 552.730 4.280 ;
        RECT 553.570 3.670 555.030 4.280 ;
        RECT 555.870 3.670 557.330 4.280 ;
        RECT 558.170 3.670 559.630 4.280 ;
        RECT 560.470 3.670 561.930 4.280 ;
        RECT 562.770 3.670 564.230 4.280 ;
        RECT 565.070 3.670 566.530 4.280 ;
        RECT 567.370 3.670 568.830 4.280 ;
        RECT 569.670 3.670 571.130 4.280 ;
        RECT 571.970 3.670 573.430 4.280 ;
        RECT 574.270 3.670 575.730 4.280 ;
        RECT 576.570 3.670 578.030 4.280 ;
        RECT 578.870 3.670 580.330 4.280 ;
        RECT 581.170 3.670 582.630 4.280 ;
        RECT 583.470 3.670 584.930 4.280 ;
        RECT 585.770 3.670 587.230 4.280 ;
        RECT 588.070 3.670 589.530 4.280 ;
        RECT 590.370 3.670 591.830 4.280 ;
        RECT 592.670 3.670 594.130 4.280 ;
        RECT 594.970 3.670 596.430 4.280 ;
        RECT 597.270 3.670 598.730 4.280 ;
        RECT 599.570 3.670 601.030 4.280 ;
        RECT 601.870 3.670 603.330 4.280 ;
        RECT 604.170 3.670 605.630 4.280 ;
        RECT 606.470 3.670 607.930 4.280 ;
        RECT 608.770 3.670 610.230 4.280 ;
        RECT 611.070 3.670 612.530 4.280 ;
        RECT 613.370 3.670 614.830 4.280 ;
        RECT 615.670 3.670 617.130 4.280 ;
        RECT 617.970 3.670 619.430 4.280 ;
        RECT 620.270 3.670 621.730 4.280 ;
        RECT 622.570 3.670 624.030 4.280 ;
        RECT 624.870 3.670 626.330 4.280 ;
        RECT 627.170 3.670 628.630 4.280 ;
        RECT 629.470 3.670 630.930 4.280 ;
        RECT 631.770 3.670 633.230 4.280 ;
        RECT 634.070 3.670 635.530 4.280 ;
        RECT 636.370 3.670 637.830 4.280 ;
        RECT 638.670 3.670 640.130 4.280 ;
        RECT 640.970 3.670 642.430 4.280 ;
        RECT 643.270 3.670 644.730 4.280 ;
        RECT 645.570 3.670 647.030 4.280 ;
        RECT 647.870 3.670 649.330 4.280 ;
        RECT 650.170 3.670 651.630 4.280 ;
        RECT 652.470 3.670 653.930 4.280 ;
        RECT 654.770 3.670 656.230 4.280 ;
        RECT 657.070 3.670 658.530 4.280 ;
        RECT 659.370 3.670 660.830 4.280 ;
        RECT 661.670 3.670 663.130 4.280 ;
        RECT 663.970 3.670 665.430 4.280 ;
        RECT 666.270 3.670 667.730 4.280 ;
        RECT 668.570 3.670 670.030 4.280 ;
        RECT 670.870 3.670 672.330 4.280 ;
        RECT 673.170 3.670 674.630 4.280 ;
        RECT 675.470 3.670 676.930 4.280 ;
        RECT 677.770 3.670 679.230 4.280 ;
        RECT 680.070 3.670 681.530 4.280 ;
        RECT 682.370 3.670 683.830 4.280 ;
        RECT 684.670 3.670 686.130 4.280 ;
        RECT 686.970 3.670 688.430 4.280 ;
        RECT 689.270 3.670 690.730 4.280 ;
        RECT 691.570 3.670 693.030 4.280 ;
        RECT 693.870 3.670 695.330 4.280 ;
        RECT 696.170 3.670 697.630 4.280 ;
        RECT 698.470 3.670 699.930 4.280 ;
        RECT 700.770 3.670 702.230 4.280 ;
        RECT 703.070 3.670 704.530 4.280 ;
        RECT 705.370 3.670 706.830 4.280 ;
        RECT 707.670 3.670 709.130 4.280 ;
        RECT 709.970 3.670 711.430 4.280 ;
        RECT 712.270 3.670 713.730 4.280 ;
        RECT 714.570 3.670 716.030 4.280 ;
        RECT 716.870 3.670 718.330 4.280 ;
        RECT 719.170 3.670 720.630 4.280 ;
        RECT 721.470 3.670 722.930 4.280 ;
        RECT 723.770 3.670 725.230 4.280 ;
        RECT 726.070 3.670 727.530 4.280 ;
        RECT 728.370 3.670 729.830 4.280 ;
        RECT 730.670 3.670 732.130 4.280 ;
        RECT 732.970 3.670 734.430 4.280 ;
        RECT 735.270 3.670 736.730 4.280 ;
        RECT 737.570 3.670 739.030 4.280 ;
        RECT 739.870 3.670 741.330 4.280 ;
        RECT 742.170 3.670 743.630 4.280 ;
        RECT 744.470 3.670 745.930 4.280 ;
        RECT 746.770 3.670 748.230 4.280 ;
        RECT 749.070 3.670 750.530 4.280 ;
        RECT 751.370 3.670 752.830 4.280 ;
        RECT 753.670 3.670 755.130 4.280 ;
        RECT 755.970 3.670 757.430 4.280 ;
        RECT 758.270 3.670 759.730 4.280 ;
        RECT 760.570 3.670 762.030 4.280 ;
        RECT 762.870 3.670 764.330 4.280 ;
        RECT 765.170 3.670 766.630 4.280 ;
        RECT 767.470 3.670 768.930 4.280 ;
        RECT 769.770 3.670 771.230 4.280 ;
        RECT 772.070 3.670 773.530 4.280 ;
        RECT 774.370 3.670 775.830 4.280 ;
        RECT 776.670 3.670 778.130 4.280 ;
        RECT 778.970 3.670 780.430 4.280 ;
        RECT 781.270 3.670 782.730 4.280 ;
        RECT 783.570 3.670 785.030 4.280 ;
        RECT 785.870 3.670 787.330 4.280 ;
        RECT 788.170 3.670 789.630 4.280 ;
        RECT 790.470 3.670 791.930 4.280 ;
        RECT 792.770 3.670 794.230 4.280 ;
        RECT 795.070 3.670 796.530 4.280 ;
        RECT 797.370 3.670 798.830 4.280 ;
        RECT 799.670 3.670 801.130 4.280 ;
        RECT 801.970 3.670 803.430 4.280 ;
        RECT 804.270 3.670 805.730 4.280 ;
        RECT 806.570 3.670 808.030 4.280 ;
        RECT 808.870 3.670 810.330 4.280 ;
        RECT 811.170 3.670 812.630 4.280 ;
        RECT 813.470 3.670 814.930 4.280 ;
        RECT 815.770 3.670 817.230 4.280 ;
        RECT 818.070 3.670 819.530 4.280 ;
        RECT 820.370 3.670 821.830 4.280 ;
        RECT 822.670 3.670 824.130 4.280 ;
        RECT 824.970 3.670 826.430 4.280 ;
        RECT 827.270 3.670 828.730 4.280 ;
        RECT 829.570 3.670 831.030 4.280 ;
        RECT 831.870 3.670 833.330 4.280 ;
        RECT 834.170 3.670 835.630 4.280 ;
        RECT 836.470 3.670 837.930 4.280 ;
        RECT 838.770 3.670 840.230 4.280 ;
        RECT 841.070 3.670 842.530 4.280 ;
        RECT 843.370 3.670 844.830 4.280 ;
        RECT 845.670 3.670 847.130 4.280 ;
        RECT 847.970 3.670 849.430 4.280 ;
        RECT 850.270 3.670 851.730 4.280 ;
        RECT 852.570 3.670 854.030 4.280 ;
        RECT 854.870 3.670 856.330 4.280 ;
        RECT 857.170 3.670 858.630 4.280 ;
        RECT 859.470 3.670 860.930 4.280 ;
        RECT 861.770 3.670 863.230 4.280 ;
        RECT 864.070 3.670 865.530 4.280 ;
        RECT 866.370 3.670 867.830 4.280 ;
        RECT 868.670 3.670 870.130 4.280 ;
        RECT 870.970 3.670 872.430 4.280 ;
        RECT 873.270 3.670 874.730 4.280 ;
        RECT 875.570 3.670 877.030 4.280 ;
        RECT 877.870 3.670 879.330 4.280 ;
        RECT 880.170 3.670 881.630 4.280 ;
        RECT 882.470 3.670 883.930 4.280 ;
        RECT 884.770 3.670 886.230 4.280 ;
        RECT 887.070 3.670 888.530 4.280 ;
        RECT 889.370 3.670 890.830 4.280 ;
        RECT 891.670 3.670 893.130 4.280 ;
        RECT 893.970 3.670 895.430 4.280 ;
        RECT 896.270 3.670 897.730 4.280 ;
        RECT 898.570 3.670 900.030 4.280 ;
        RECT 900.870 3.670 902.330 4.280 ;
        RECT 903.170 3.670 904.630 4.280 ;
        RECT 905.470 3.670 906.930 4.280 ;
        RECT 907.770 3.670 909.230 4.280 ;
        RECT 910.070 3.670 911.530 4.280 ;
        RECT 912.370 3.670 913.830 4.280 ;
        RECT 914.670 3.670 916.130 4.280 ;
        RECT 916.970 3.670 918.430 4.280 ;
        RECT 919.270 3.670 920.730 4.280 ;
        RECT 921.570 3.670 923.030 4.280 ;
        RECT 923.870 3.670 925.330 4.280 ;
        RECT 926.170 3.670 927.630 4.280 ;
        RECT 928.470 3.670 929.930 4.280 ;
        RECT 930.770 3.670 932.230 4.280 ;
        RECT 933.070 3.670 934.530 4.280 ;
        RECT 935.370 3.670 936.830 4.280 ;
        RECT 937.670 3.670 939.130 4.280 ;
        RECT 939.970 3.670 941.430 4.280 ;
        RECT 942.270 3.670 943.730 4.280 ;
        RECT 944.570 3.670 946.030 4.280 ;
        RECT 946.870 3.670 948.330 4.280 ;
        RECT 949.170 3.670 950.630 4.280 ;
        RECT 951.470 3.670 952.930 4.280 ;
        RECT 953.770 3.670 955.230 4.280 ;
        RECT 956.070 3.670 957.530 4.280 ;
        RECT 958.370 3.670 959.830 4.280 ;
        RECT 960.670 3.670 962.130 4.280 ;
        RECT 962.970 3.670 964.430 4.280 ;
        RECT 965.270 3.670 966.730 4.280 ;
        RECT 967.570 3.670 969.030 4.280 ;
        RECT 969.870 3.670 971.330 4.280 ;
        RECT 972.170 3.670 973.630 4.280 ;
        RECT 974.470 3.670 975.930 4.280 ;
        RECT 976.770 3.670 978.230 4.280 ;
        RECT 979.070 3.670 980.530 4.280 ;
        RECT 981.370 3.670 982.830 4.280 ;
        RECT 983.670 3.670 985.130 4.280 ;
        RECT 985.970 3.670 987.430 4.280 ;
        RECT 988.270 3.670 989.730 4.280 ;
        RECT 990.570 3.670 992.030 4.280 ;
        RECT 992.870 3.670 994.330 4.280 ;
        RECT 995.170 3.670 996.630 4.280 ;
        RECT 997.470 3.670 998.930 4.280 ;
        RECT 999.770 3.670 1001.230 4.280 ;
        RECT 1002.070 3.670 1003.530 4.280 ;
        RECT 1004.370 3.670 1005.830 4.280 ;
        RECT 1006.670 3.670 1008.130 4.280 ;
        RECT 1008.970 3.670 1010.430 4.280 ;
        RECT 1011.270 3.670 1012.730 4.280 ;
        RECT 1013.570 3.670 1015.030 4.280 ;
        RECT 1015.870 3.670 1017.330 4.280 ;
        RECT 1018.170 3.670 1019.630 4.280 ;
        RECT 1020.470 3.670 1021.930 4.280 ;
        RECT 1022.770 3.670 1024.230 4.280 ;
        RECT 1025.070 3.670 1026.530 4.280 ;
        RECT 1027.370 3.670 1028.830 4.280 ;
        RECT 1029.670 3.670 1031.130 4.280 ;
        RECT 1031.970 3.670 1033.430 4.280 ;
        RECT 1034.270 3.670 1035.730 4.280 ;
        RECT 1036.570 3.670 1038.030 4.280 ;
        RECT 1038.870 3.670 1040.330 4.280 ;
        RECT 1041.170 3.670 1042.630 4.280 ;
        RECT 1043.470 3.670 1044.930 4.280 ;
        RECT 1045.770 3.670 1047.230 4.280 ;
        RECT 1048.070 3.670 1049.530 4.280 ;
        RECT 1050.370 3.670 1051.830 4.280 ;
        RECT 1052.670 3.670 1054.130 4.280 ;
        RECT 1054.970 3.670 1056.430 4.280 ;
        RECT 1057.270 3.670 1058.730 4.280 ;
        RECT 1059.570 3.670 1061.030 4.280 ;
        RECT 1061.870 3.670 1063.330 4.280 ;
        RECT 1064.170 3.670 1065.630 4.280 ;
        RECT 1066.470 3.670 1067.930 4.280 ;
        RECT 1068.770 3.670 1070.230 4.280 ;
        RECT 1071.070 3.670 1072.530 4.280 ;
        RECT 1073.370 3.670 1074.830 4.280 ;
        RECT 1075.670 3.670 1077.130 4.280 ;
        RECT 1077.970 3.670 1079.430 4.280 ;
        RECT 1080.270 3.670 1081.730 4.280 ;
        RECT 1082.570 3.670 1084.030 4.280 ;
        RECT 1084.870 3.670 1086.330 4.280 ;
        RECT 1087.170 3.670 1088.630 4.280 ;
        RECT 1089.470 3.670 1090.930 4.280 ;
        RECT 1091.770 3.670 1093.230 4.280 ;
        RECT 1094.070 3.670 1095.530 4.280 ;
        RECT 1096.370 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1100.130 4.280 ;
        RECT 1100.970 3.670 1102.430 4.280 ;
        RECT 1103.270 3.670 1104.730 4.280 ;
        RECT 1105.570 3.670 1107.030 4.280 ;
        RECT 1107.870 3.670 1109.330 4.280 ;
        RECT 1110.170 3.670 1111.630 4.280 ;
        RECT 1112.470 3.670 1113.930 4.280 ;
        RECT 1114.770 3.670 1116.230 4.280 ;
        RECT 1117.070 3.670 1118.530 4.280 ;
        RECT 1119.370 3.670 1120.830 4.280 ;
        RECT 1121.670 3.670 1123.130 4.280 ;
        RECT 1123.970 3.670 1125.430 4.280 ;
        RECT 1126.270 3.670 1127.730 4.280 ;
        RECT 1128.570 3.670 1130.030 4.280 ;
        RECT 1130.870 3.670 1132.330 4.280 ;
        RECT 1133.170 3.670 1134.630 4.280 ;
        RECT 1135.470 3.670 1136.930 4.280 ;
        RECT 1137.770 3.670 1139.230 4.280 ;
        RECT 1140.070 3.670 1141.530 4.280 ;
        RECT 1142.370 3.670 1143.830 4.280 ;
        RECT 1144.670 3.670 1146.130 4.280 ;
        RECT 1146.970 3.670 1148.430 4.280 ;
        RECT 1149.270 3.670 1150.730 4.280 ;
        RECT 1151.570 3.670 1153.030 4.280 ;
        RECT 1153.870 3.670 1155.330 4.280 ;
        RECT 1156.170 3.670 1157.630 4.280 ;
        RECT 1158.470 3.670 1159.930 4.280 ;
        RECT 1160.770 3.670 1162.230 4.280 ;
        RECT 1163.070 3.670 1164.530 4.280 ;
        RECT 1165.370 3.670 1166.830 4.280 ;
        RECT 1167.670 3.670 1169.130 4.280 ;
        RECT 1169.970 3.670 1171.430 4.280 ;
        RECT 1172.270 3.670 1173.730 4.280 ;
        RECT 1174.570 3.670 1176.030 4.280 ;
        RECT 1176.870 3.670 1178.330 4.280 ;
        RECT 1179.170 3.670 1180.630 4.280 ;
        RECT 1181.470 3.670 1182.930 4.280 ;
        RECT 1183.770 3.670 1185.230 4.280 ;
        RECT 1186.070 3.670 1187.530 4.280 ;
        RECT 1188.370 3.670 1189.830 4.280 ;
        RECT 1190.670 3.670 1192.130 4.280 ;
        RECT 1192.970 3.670 1194.430 4.280 ;
        RECT 1195.270 3.670 1196.730 4.280 ;
        RECT 1197.570 3.670 1199.030 4.280 ;
        RECT 1199.870 3.670 1201.330 4.280 ;
        RECT 1202.170 3.670 1203.630 4.280 ;
        RECT 1204.470 3.670 1205.930 4.280 ;
        RECT 1206.770 3.670 1208.230 4.280 ;
        RECT 1209.070 3.670 1210.530 4.280 ;
        RECT 1211.370 3.670 1212.830 4.280 ;
        RECT 1213.670 3.670 1215.130 4.280 ;
        RECT 1215.970 3.670 1273.640 4.280 ;
      LAYER met3 ;
        RECT 11.565 10.715 1251.430 1387.365 ;
      LAYER met4 ;
        RECT 15.935 11.055 20.640 1385.665 ;
        RECT 23.040 11.055 97.440 1385.665 ;
        RECT 99.840 11.055 174.240 1385.665 ;
        RECT 176.640 11.055 251.040 1385.665 ;
        RECT 253.440 11.055 327.840 1385.665 ;
        RECT 330.240 11.055 404.640 1385.665 ;
        RECT 407.040 11.055 481.440 1385.665 ;
        RECT 483.840 11.055 558.240 1385.665 ;
        RECT 560.640 11.055 635.040 1385.665 ;
        RECT 637.440 11.055 711.840 1385.665 ;
        RECT 714.240 11.055 788.640 1385.665 ;
        RECT 791.040 11.055 865.440 1385.665 ;
        RECT 867.840 11.055 942.240 1385.665 ;
        RECT 944.640 11.055 1019.040 1385.665 ;
        RECT 1021.440 11.055 1095.840 1385.665 ;
        RECT 1098.240 11.055 1119.345 1385.665 ;
  END
END wb_pio
END LIBRARY

