magic
tech sky130B
magscale 1 2
timestamp 1672205199
<< nwell >>
rect 1066 276613 258926 277179
rect 1066 275525 258926 276091
rect 1066 274437 258926 275003
rect 1066 273349 258926 273915
rect 1066 272261 258926 272827
rect 1066 271173 258926 271739
rect 1066 270085 258926 270651
rect 1066 268997 258926 269563
rect 1066 267909 258926 268475
rect 1066 266821 258926 267387
rect 1066 265733 258926 266299
rect 1066 264645 258926 265211
rect 1066 263557 258926 264123
rect 1066 262469 258926 263035
rect 1066 261381 258926 261947
rect 1066 260293 258926 260859
rect 1066 259205 258926 259771
rect 1066 258117 258926 258683
rect 1066 257029 258926 257595
rect 1066 255941 258926 256507
rect 1066 254853 258926 255419
rect 1066 253765 258926 254331
rect 1066 252677 258926 253243
rect 1066 251589 258926 252155
rect 1066 250501 258926 251067
rect 1066 249413 258926 249979
rect 1066 248325 258926 248891
rect 1066 247237 258926 247803
rect 1066 246149 258926 246715
rect 1066 245061 258926 245627
rect 1066 243973 258926 244539
rect 1066 242885 258926 243451
rect 1066 241797 258926 242363
rect 1066 240709 258926 241275
rect 1066 239621 258926 240187
rect 1066 238533 258926 239099
rect 1066 237445 258926 238011
rect 1066 236357 258926 236923
rect 1066 235269 258926 235835
rect 1066 234181 258926 234747
rect 1066 233093 258926 233659
rect 1066 232005 258926 232571
rect 1066 230917 258926 231483
rect 1066 229829 258926 230395
rect 1066 228741 258926 229307
rect 1066 227653 258926 228219
rect 1066 226565 258926 227131
rect 1066 225477 258926 226043
rect 1066 224389 258926 224955
rect 1066 223301 258926 223867
rect 1066 222213 258926 222779
rect 1066 221125 258926 221691
rect 1066 220037 258926 220603
rect 1066 218949 258926 219515
rect 1066 217861 258926 218427
rect 1066 216773 258926 217339
rect 1066 215685 258926 216251
rect 1066 214597 258926 215163
rect 1066 213509 258926 214075
rect 1066 212421 258926 212987
rect 1066 211333 258926 211899
rect 1066 210245 258926 210811
rect 1066 209157 258926 209723
rect 1066 208069 258926 208635
rect 1066 206981 258926 207547
rect 1066 205893 258926 206459
rect 1066 204805 258926 205371
rect 1066 203717 258926 204283
rect 1066 202629 258926 203195
rect 1066 201541 258926 202107
rect 1066 200453 258926 201019
rect 1066 199365 258926 199931
rect 1066 198277 258926 198843
rect 1066 197189 258926 197755
rect 1066 196101 258926 196667
rect 1066 195013 258926 195579
rect 1066 193925 258926 194491
rect 1066 192837 258926 193403
rect 1066 191749 258926 192315
rect 1066 190661 258926 191227
rect 1066 189573 258926 190139
rect 1066 188485 258926 189051
rect 1066 187397 258926 187963
rect 1066 186309 258926 186875
rect 1066 185221 258926 185787
rect 1066 184133 258926 184699
rect 1066 183045 258926 183611
rect 1066 181957 258926 182523
rect 1066 180869 258926 181435
rect 1066 179781 258926 180347
rect 1066 178693 258926 179259
rect 1066 177605 258926 178171
rect 1066 176517 258926 177083
rect 1066 175429 258926 175995
rect 1066 174341 258926 174907
rect 1066 173253 258926 173819
rect 1066 172165 258926 172731
rect 1066 171077 258926 171643
rect 1066 169989 258926 170555
rect 1066 168901 258926 169467
rect 1066 167813 258926 168379
rect 1066 166725 258926 167291
rect 1066 165637 258926 166203
rect 1066 164549 258926 165115
rect 1066 163461 258926 164027
rect 1066 162373 258926 162939
rect 1066 161285 258926 161851
rect 1066 160197 258926 160763
rect 1066 159109 258926 159675
rect 1066 158021 258926 158587
rect 1066 156933 258926 157499
rect 1066 155845 258926 156411
rect 1066 154757 258926 155323
rect 1066 153669 258926 154235
rect 1066 152581 258926 153147
rect 1066 151493 258926 152059
rect 1066 150405 258926 150971
rect 1066 149317 258926 149883
rect 1066 148229 258926 148795
rect 1066 147141 258926 147707
rect 1066 146053 258926 146619
rect 1066 144965 258926 145531
rect 1066 143877 258926 144443
rect 1066 142789 258926 143355
rect 1066 141701 258926 142267
rect 1066 140613 258926 141179
rect 1066 139525 258926 140091
rect 1066 138437 258926 139003
rect 1066 137349 258926 137915
rect 1066 136261 258926 136827
rect 1066 135173 258926 135739
rect 1066 134085 258926 134651
rect 1066 132997 258926 133563
rect 1066 131909 258926 132475
rect 1066 130821 258926 131387
rect 1066 129733 258926 130299
rect 1066 128645 258926 129211
rect 1066 127557 258926 128123
rect 1066 126469 258926 127035
rect 1066 125381 258926 125947
rect 1066 124293 258926 124859
rect 1066 123205 258926 123771
rect 1066 122117 258926 122683
rect 1066 121029 258926 121595
rect 1066 119941 258926 120507
rect 1066 118853 258926 119419
rect 1066 117765 258926 118331
rect 1066 116677 258926 117243
rect 1066 115589 258926 116155
rect 1066 114501 258926 115067
rect 1066 113413 258926 113979
rect 1066 112325 258926 112891
rect 1066 111237 258926 111803
rect 1066 110149 258926 110715
rect 1066 109061 258926 109627
rect 1066 107973 258926 108539
rect 1066 106885 258926 107451
rect 1066 105797 258926 106363
rect 1066 104709 258926 105275
rect 1066 103621 258926 104187
rect 1066 102533 258926 103099
rect 1066 101445 258926 102011
rect 1066 100357 258926 100923
rect 1066 99269 258926 99835
rect 1066 98181 258926 98747
rect 1066 97093 258926 97659
rect 1066 96005 258926 96571
rect 1066 94917 258926 95483
rect 1066 93829 258926 94395
rect 1066 92741 258926 93307
rect 1066 91653 258926 92219
rect 1066 90565 258926 91131
rect 1066 89477 258926 90043
rect 1066 88389 258926 88955
rect 1066 87301 258926 87867
rect 1066 86213 258926 86779
rect 1066 85125 258926 85691
rect 1066 84037 258926 84603
rect 1066 82949 258926 83515
rect 1066 81861 258926 82427
rect 1066 80773 258926 81339
rect 1066 79685 258926 80251
rect 1066 78597 258926 79163
rect 1066 77509 258926 78075
rect 1066 76421 258926 76987
rect 1066 75333 258926 75899
rect 1066 74245 258926 74811
rect 1066 73157 258926 73723
rect 1066 72069 258926 72635
rect 1066 70981 258926 71547
rect 1066 69893 258926 70459
rect 1066 68805 258926 69371
rect 1066 67717 258926 68283
rect 1066 66629 258926 67195
rect 1066 65541 258926 66107
rect 1066 64453 258926 65019
rect 1066 63365 258926 63931
rect 1066 62277 258926 62843
rect 1066 61189 258926 61755
rect 1066 60101 258926 60667
rect 1066 59013 258926 59579
rect 1066 57925 258926 58491
rect 1066 56837 258926 57403
rect 1066 55749 258926 56315
rect 1066 54661 258926 55227
rect 1066 53573 258926 54139
rect 1066 52485 258926 53051
rect 1066 51397 258926 51963
rect 1066 50309 258926 50875
rect 1066 49221 258926 49787
rect 1066 48133 258926 48699
rect 1066 47045 258926 47611
rect 1066 45957 258926 46523
rect 1066 44869 258926 45435
rect 1066 43781 258926 44347
rect 1066 42693 258926 43259
rect 1066 41605 258926 42171
rect 1066 40517 258926 41083
rect 1066 39429 258926 39995
rect 1066 38341 258926 38907
rect 1066 37253 258926 37819
rect 1066 36165 258926 36731
rect 1066 35077 258926 35643
rect 1066 33989 258926 34555
rect 1066 32901 258926 33467
rect 1066 31813 258926 32379
rect 1066 30725 258926 31291
rect 1066 29637 258926 30203
rect 1066 28549 258926 29115
rect 1066 27461 258926 28027
rect 1066 26373 258926 26939
rect 1066 25285 258926 25851
rect 1066 24197 258926 24763
rect 1066 23109 258926 23675
rect 1066 22021 258926 22587
rect 1066 20933 258926 21499
rect 1066 19845 258926 20411
rect 1066 18757 258926 19323
rect 1066 17669 258926 18235
rect 1066 16581 258926 17147
rect 1066 15493 258926 16059
rect 1066 14405 258926 14971
rect 1066 13317 258926 13883
rect 1066 12229 258926 12795
rect 1066 11141 258926 11707
rect 1066 10053 258926 10619
rect 1066 8965 258926 9531
rect 1066 7877 258926 8443
rect 1066 6789 258926 7355
rect 1066 5701 258926 6267
rect 1066 4613 258926 5179
rect 1066 3525 258926 4091
rect 1066 2437 258926 3003
<< obsli1 >>
rect 1104 2159 258888 277457
<< obsm1 >>
rect 1104 1640 258888 277488
<< metal2 >>
rect 5170 279200 5226 280000
rect 7378 279200 7434 280000
rect 9586 279200 9642 280000
rect 11794 279200 11850 280000
rect 14002 279200 14058 280000
rect 16210 279200 16266 280000
rect 18418 279200 18474 280000
rect 20626 279200 20682 280000
rect 22834 279200 22890 280000
rect 25042 279200 25098 280000
rect 27250 279200 27306 280000
rect 29458 279200 29514 280000
rect 31666 279200 31722 280000
rect 33874 279200 33930 280000
rect 36082 279200 36138 280000
rect 38290 279200 38346 280000
rect 40498 279200 40554 280000
rect 42706 279200 42762 280000
rect 44914 279200 44970 280000
rect 47122 279200 47178 280000
rect 49330 279200 49386 280000
rect 51538 279200 51594 280000
rect 53746 279200 53802 280000
rect 55954 279200 56010 280000
rect 58162 279200 58218 280000
rect 60370 279200 60426 280000
rect 62578 279200 62634 280000
rect 64786 279200 64842 280000
rect 66994 279200 67050 280000
rect 69202 279200 69258 280000
rect 71410 279200 71466 280000
rect 73618 279200 73674 280000
rect 75826 279200 75882 280000
rect 78034 279200 78090 280000
rect 80242 279200 80298 280000
rect 82450 279200 82506 280000
rect 84658 279200 84714 280000
rect 86866 279200 86922 280000
rect 89074 279200 89130 280000
rect 91282 279200 91338 280000
rect 93490 279200 93546 280000
rect 95698 279200 95754 280000
rect 97906 279200 97962 280000
rect 100114 279200 100170 280000
rect 102322 279200 102378 280000
rect 104530 279200 104586 280000
rect 106738 279200 106794 280000
rect 108946 279200 109002 280000
rect 111154 279200 111210 280000
rect 113362 279200 113418 280000
rect 115570 279200 115626 280000
rect 117778 279200 117834 280000
rect 119986 279200 120042 280000
rect 122194 279200 122250 280000
rect 124402 279200 124458 280000
rect 126610 279200 126666 280000
rect 128818 279200 128874 280000
rect 131026 279200 131082 280000
rect 133234 279200 133290 280000
rect 135442 279200 135498 280000
rect 137650 279200 137706 280000
rect 139858 279200 139914 280000
rect 142066 279200 142122 280000
rect 144274 279200 144330 280000
rect 146482 279200 146538 280000
rect 148690 279200 148746 280000
rect 150898 279200 150954 280000
rect 153106 279200 153162 280000
rect 155314 279200 155370 280000
rect 157522 279200 157578 280000
rect 159730 279200 159786 280000
rect 161938 279200 161994 280000
rect 164146 279200 164202 280000
rect 166354 279200 166410 280000
rect 168562 279200 168618 280000
rect 170770 279200 170826 280000
rect 172978 279200 173034 280000
rect 175186 279200 175242 280000
rect 177394 279200 177450 280000
rect 179602 279200 179658 280000
rect 181810 279200 181866 280000
rect 184018 279200 184074 280000
rect 186226 279200 186282 280000
rect 188434 279200 188490 280000
rect 190642 279200 190698 280000
rect 192850 279200 192906 280000
rect 195058 279200 195114 280000
rect 197266 279200 197322 280000
rect 199474 279200 199530 280000
rect 201682 279200 201738 280000
rect 203890 279200 203946 280000
rect 206098 279200 206154 280000
rect 208306 279200 208362 280000
rect 210514 279200 210570 280000
rect 212722 279200 212778 280000
rect 214930 279200 214986 280000
rect 217138 279200 217194 280000
rect 219346 279200 219402 280000
rect 221554 279200 221610 280000
rect 223762 279200 223818 280000
rect 225970 279200 226026 280000
rect 228178 279200 228234 280000
rect 230386 279200 230442 280000
rect 232594 279200 232650 280000
rect 234802 279200 234858 280000
rect 237010 279200 237066 280000
rect 239218 279200 239274 280000
rect 241426 279200 241482 280000
rect 243634 279200 243690 280000
rect 245842 279200 245898 280000
rect 248050 279200 248106 280000
rect 250258 279200 250314 280000
rect 252466 279200 252522 280000
rect 254674 279200 254730 280000
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
rect 23202 0 23258 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25502 0 25558 800
rect 25962 0 26018 800
rect 26422 0 26478 800
rect 26882 0 26938 800
rect 27342 0 27398 800
rect 27802 0 27858 800
rect 28262 0 28318 800
rect 28722 0 28778 800
rect 29182 0 29238 800
rect 29642 0 29698 800
rect 30102 0 30158 800
rect 30562 0 30618 800
rect 31022 0 31078 800
rect 31482 0 31538 800
rect 31942 0 31998 800
rect 32402 0 32458 800
rect 32862 0 32918 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34242 0 34298 800
rect 34702 0 34758 800
rect 35162 0 35218 800
rect 35622 0 35678 800
rect 36082 0 36138 800
rect 36542 0 36598 800
rect 37002 0 37058 800
rect 37462 0 37518 800
rect 37922 0 37978 800
rect 38382 0 38438 800
rect 38842 0 38898 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40682 0 40738 800
rect 41142 0 41198 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42522 0 42578 800
rect 42982 0 43038 800
rect 43442 0 43498 800
rect 43902 0 43958 800
rect 44362 0 44418 800
rect 44822 0 44878 800
rect 45282 0 45338 800
rect 45742 0 45798 800
rect 46202 0 46258 800
rect 46662 0 46718 800
rect 47122 0 47178 800
rect 47582 0 47638 800
rect 48042 0 48098 800
rect 48502 0 48558 800
rect 48962 0 49018 800
rect 49422 0 49478 800
rect 49882 0 49938 800
rect 50342 0 50398 800
rect 50802 0 50858 800
rect 51262 0 51318 800
rect 51722 0 51778 800
rect 52182 0 52238 800
rect 52642 0 52698 800
rect 53102 0 53158 800
rect 53562 0 53618 800
rect 54022 0 54078 800
rect 54482 0 54538 800
rect 54942 0 54998 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56322 0 56378 800
rect 56782 0 56838 800
rect 57242 0 57298 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58622 0 58678 800
rect 59082 0 59138 800
rect 59542 0 59598 800
rect 60002 0 60058 800
rect 60462 0 60518 800
rect 60922 0 60978 800
rect 61382 0 61438 800
rect 61842 0 61898 800
rect 62302 0 62358 800
rect 62762 0 62818 800
rect 63222 0 63278 800
rect 63682 0 63738 800
rect 64142 0 64198 800
rect 64602 0 64658 800
rect 65062 0 65118 800
rect 65522 0 65578 800
rect 65982 0 66038 800
rect 66442 0 66498 800
rect 66902 0 66958 800
rect 67362 0 67418 800
rect 67822 0 67878 800
rect 68282 0 68338 800
rect 68742 0 68798 800
rect 69202 0 69258 800
rect 69662 0 69718 800
rect 70122 0 70178 800
rect 70582 0 70638 800
rect 71042 0 71098 800
rect 71502 0 71558 800
rect 71962 0 72018 800
rect 72422 0 72478 800
rect 72882 0 72938 800
rect 73342 0 73398 800
rect 73802 0 73858 800
rect 74262 0 74318 800
rect 74722 0 74778 800
rect 75182 0 75238 800
rect 75642 0 75698 800
rect 76102 0 76158 800
rect 76562 0 76618 800
rect 77022 0 77078 800
rect 77482 0 77538 800
rect 77942 0 77998 800
rect 78402 0 78458 800
rect 78862 0 78918 800
rect 79322 0 79378 800
rect 79782 0 79838 800
rect 80242 0 80298 800
rect 80702 0 80758 800
rect 81162 0 81218 800
rect 81622 0 81678 800
rect 82082 0 82138 800
rect 82542 0 82598 800
rect 83002 0 83058 800
rect 83462 0 83518 800
rect 83922 0 83978 800
rect 84382 0 84438 800
rect 84842 0 84898 800
rect 85302 0 85358 800
rect 85762 0 85818 800
rect 86222 0 86278 800
rect 86682 0 86738 800
rect 87142 0 87198 800
rect 87602 0 87658 800
rect 88062 0 88118 800
rect 88522 0 88578 800
rect 88982 0 89038 800
rect 89442 0 89498 800
rect 89902 0 89958 800
rect 90362 0 90418 800
rect 90822 0 90878 800
rect 91282 0 91338 800
rect 91742 0 91798 800
rect 92202 0 92258 800
rect 92662 0 92718 800
rect 93122 0 93178 800
rect 93582 0 93638 800
rect 94042 0 94098 800
rect 94502 0 94558 800
rect 94962 0 95018 800
rect 95422 0 95478 800
rect 95882 0 95938 800
rect 96342 0 96398 800
rect 96802 0 96858 800
rect 97262 0 97318 800
rect 97722 0 97778 800
rect 98182 0 98238 800
rect 98642 0 98698 800
rect 99102 0 99158 800
rect 99562 0 99618 800
rect 100022 0 100078 800
rect 100482 0 100538 800
rect 100942 0 100998 800
rect 101402 0 101458 800
rect 101862 0 101918 800
rect 102322 0 102378 800
rect 102782 0 102838 800
rect 103242 0 103298 800
rect 103702 0 103758 800
rect 104162 0 104218 800
rect 104622 0 104678 800
rect 105082 0 105138 800
rect 105542 0 105598 800
rect 106002 0 106058 800
rect 106462 0 106518 800
rect 106922 0 106978 800
rect 107382 0 107438 800
rect 107842 0 107898 800
rect 108302 0 108358 800
rect 108762 0 108818 800
rect 109222 0 109278 800
rect 109682 0 109738 800
rect 110142 0 110198 800
rect 110602 0 110658 800
rect 111062 0 111118 800
rect 111522 0 111578 800
rect 111982 0 112038 800
rect 112442 0 112498 800
rect 112902 0 112958 800
rect 113362 0 113418 800
rect 113822 0 113878 800
rect 114282 0 114338 800
rect 114742 0 114798 800
rect 115202 0 115258 800
rect 115662 0 115718 800
rect 116122 0 116178 800
rect 116582 0 116638 800
rect 117042 0 117098 800
rect 117502 0 117558 800
rect 117962 0 118018 800
rect 118422 0 118478 800
rect 118882 0 118938 800
rect 119342 0 119398 800
rect 119802 0 119858 800
rect 120262 0 120318 800
rect 120722 0 120778 800
rect 121182 0 121238 800
rect 121642 0 121698 800
rect 122102 0 122158 800
rect 122562 0 122618 800
rect 123022 0 123078 800
rect 123482 0 123538 800
rect 123942 0 123998 800
rect 124402 0 124458 800
rect 124862 0 124918 800
rect 125322 0 125378 800
rect 125782 0 125838 800
rect 126242 0 126298 800
rect 126702 0 126758 800
rect 127162 0 127218 800
rect 127622 0 127678 800
rect 128082 0 128138 800
rect 128542 0 128598 800
rect 129002 0 129058 800
rect 129462 0 129518 800
rect 129922 0 129978 800
rect 130382 0 130438 800
rect 130842 0 130898 800
rect 131302 0 131358 800
rect 131762 0 131818 800
rect 132222 0 132278 800
rect 132682 0 132738 800
rect 133142 0 133198 800
rect 133602 0 133658 800
rect 134062 0 134118 800
rect 134522 0 134578 800
rect 134982 0 135038 800
rect 135442 0 135498 800
rect 135902 0 135958 800
rect 136362 0 136418 800
rect 136822 0 136878 800
rect 137282 0 137338 800
rect 137742 0 137798 800
rect 138202 0 138258 800
rect 138662 0 138718 800
rect 139122 0 139178 800
rect 139582 0 139638 800
rect 140042 0 140098 800
rect 140502 0 140558 800
rect 140962 0 141018 800
rect 141422 0 141478 800
rect 141882 0 141938 800
rect 142342 0 142398 800
rect 142802 0 142858 800
rect 143262 0 143318 800
rect 143722 0 143778 800
rect 144182 0 144238 800
rect 144642 0 144698 800
rect 145102 0 145158 800
rect 145562 0 145618 800
rect 146022 0 146078 800
rect 146482 0 146538 800
rect 146942 0 146998 800
rect 147402 0 147458 800
rect 147862 0 147918 800
rect 148322 0 148378 800
rect 148782 0 148838 800
rect 149242 0 149298 800
rect 149702 0 149758 800
rect 150162 0 150218 800
rect 150622 0 150678 800
rect 151082 0 151138 800
rect 151542 0 151598 800
rect 152002 0 152058 800
rect 152462 0 152518 800
rect 152922 0 152978 800
rect 153382 0 153438 800
rect 153842 0 153898 800
rect 154302 0 154358 800
rect 154762 0 154818 800
rect 155222 0 155278 800
rect 155682 0 155738 800
rect 156142 0 156198 800
rect 156602 0 156658 800
rect 157062 0 157118 800
rect 157522 0 157578 800
rect 157982 0 158038 800
rect 158442 0 158498 800
rect 158902 0 158958 800
rect 159362 0 159418 800
rect 159822 0 159878 800
rect 160282 0 160338 800
rect 160742 0 160798 800
rect 161202 0 161258 800
rect 161662 0 161718 800
rect 162122 0 162178 800
rect 162582 0 162638 800
rect 163042 0 163098 800
rect 163502 0 163558 800
rect 163962 0 164018 800
rect 164422 0 164478 800
rect 164882 0 164938 800
rect 165342 0 165398 800
rect 165802 0 165858 800
rect 166262 0 166318 800
rect 166722 0 166778 800
rect 167182 0 167238 800
rect 167642 0 167698 800
rect 168102 0 168158 800
rect 168562 0 168618 800
rect 169022 0 169078 800
rect 169482 0 169538 800
rect 169942 0 169998 800
rect 170402 0 170458 800
rect 170862 0 170918 800
rect 171322 0 171378 800
rect 171782 0 171838 800
rect 172242 0 172298 800
rect 172702 0 172758 800
rect 173162 0 173218 800
rect 173622 0 173678 800
rect 174082 0 174138 800
rect 174542 0 174598 800
rect 175002 0 175058 800
rect 175462 0 175518 800
rect 175922 0 175978 800
rect 176382 0 176438 800
rect 176842 0 176898 800
rect 177302 0 177358 800
rect 177762 0 177818 800
rect 178222 0 178278 800
rect 178682 0 178738 800
rect 179142 0 179198 800
rect 179602 0 179658 800
rect 180062 0 180118 800
rect 180522 0 180578 800
rect 180982 0 181038 800
rect 181442 0 181498 800
rect 181902 0 181958 800
rect 182362 0 182418 800
rect 182822 0 182878 800
rect 183282 0 183338 800
rect 183742 0 183798 800
rect 184202 0 184258 800
rect 184662 0 184718 800
rect 185122 0 185178 800
rect 185582 0 185638 800
rect 186042 0 186098 800
rect 186502 0 186558 800
rect 186962 0 187018 800
rect 187422 0 187478 800
rect 187882 0 187938 800
rect 188342 0 188398 800
rect 188802 0 188858 800
rect 189262 0 189318 800
rect 189722 0 189778 800
rect 190182 0 190238 800
rect 190642 0 190698 800
rect 191102 0 191158 800
rect 191562 0 191618 800
rect 192022 0 192078 800
rect 192482 0 192538 800
rect 192942 0 192998 800
rect 193402 0 193458 800
rect 193862 0 193918 800
rect 194322 0 194378 800
rect 194782 0 194838 800
rect 195242 0 195298 800
rect 195702 0 195758 800
rect 196162 0 196218 800
rect 196622 0 196678 800
rect 197082 0 197138 800
rect 197542 0 197598 800
rect 198002 0 198058 800
rect 198462 0 198518 800
rect 198922 0 198978 800
rect 199382 0 199438 800
rect 199842 0 199898 800
rect 200302 0 200358 800
rect 200762 0 200818 800
rect 201222 0 201278 800
rect 201682 0 201738 800
rect 202142 0 202198 800
rect 202602 0 202658 800
rect 203062 0 203118 800
rect 203522 0 203578 800
rect 203982 0 204038 800
rect 204442 0 204498 800
rect 204902 0 204958 800
rect 205362 0 205418 800
rect 205822 0 205878 800
rect 206282 0 206338 800
rect 206742 0 206798 800
rect 207202 0 207258 800
rect 207662 0 207718 800
rect 208122 0 208178 800
rect 208582 0 208638 800
rect 209042 0 209098 800
rect 209502 0 209558 800
rect 209962 0 210018 800
rect 210422 0 210478 800
rect 210882 0 210938 800
rect 211342 0 211398 800
rect 211802 0 211858 800
rect 212262 0 212318 800
rect 212722 0 212778 800
rect 213182 0 213238 800
rect 213642 0 213698 800
rect 214102 0 214158 800
rect 214562 0 214618 800
rect 215022 0 215078 800
rect 215482 0 215538 800
rect 215942 0 215998 800
rect 216402 0 216458 800
rect 216862 0 216918 800
rect 217322 0 217378 800
rect 217782 0 217838 800
rect 218242 0 218298 800
rect 218702 0 218758 800
rect 219162 0 219218 800
rect 219622 0 219678 800
rect 220082 0 220138 800
rect 220542 0 220598 800
rect 221002 0 221058 800
rect 221462 0 221518 800
rect 221922 0 221978 800
rect 222382 0 222438 800
rect 222842 0 222898 800
rect 223302 0 223358 800
rect 223762 0 223818 800
rect 224222 0 224278 800
rect 224682 0 224738 800
rect 225142 0 225198 800
rect 225602 0 225658 800
rect 226062 0 226118 800
rect 226522 0 226578 800
rect 226982 0 227038 800
rect 227442 0 227498 800
rect 227902 0 227958 800
rect 228362 0 228418 800
rect 228822 0 228878 800
rect 229282 0 229338 800
rect 229742 0 229798 800
rect 230202 0 230258 800
rect 230662 0 230718 800
rect 231122 0 231178 800
rect 231582 0 231638 800
rect 232042 0 232098 800
rect 232502 0 232558 800
rect 232962 0 233018 800
rect 233422 0 233478 800
rect 233882 0 233938 800
rect 234342 0 234398 800
rect 234802 0 234858 800
rect 235262 0 235318 800
rect 235722 0 235778 800
rect 236182 0 236238 800
rect 236642 0 236698 800
rect 237102 0 237158 800
rect 237562 0 237618 800
rect 238022 0 238078 800
rect 238482 0 238538 800
rect 238942 0 238998 800
rect 239402 0 239458 800
rect 239862 0 239918 800
rect 240322 0 240378 800
rect 240782 0 240838 800
rect 241242 0 241298 800
rect 241702 0 241758 800
rect 242162 0 242218 800
rect 242622 0 242678 800
rect 243082 0 243138 800
<< obsm2 >>
rect 1676 279144 5114 279290
rect 5282 279144 7322 279290
rect 7490 279144 9530 279290
rect 9698 279144 11738 279290
rect 11906 279144 13946 279290
rect 14114 279144 16154 279290
rect 16322 279144 18362 279290
rect 18530 279144 20570 279290
rect 20738 279144 22778 279290
rect 22946 279144 24986 279290
rect 25154 279144 27194 279290
rect 27362 279144 29402 279290
rect 29570 279144 31610 279290
rect 31778 279144 33818 279290
rect 33986 279144 36026 279290
rect 36194 279144 38234 279290
rect 38402 279144 40442 279290
rect 40610 279144 42650 279290
rect 42818 279144 44858 279290
rect 45026 279144 47066 279290
rect 47234 279144 49274 279290
rect 49442 279144 51482 279290
rect 51650 279144 53690 279290
rect 53858 279144 55898 279290
rect 56066 279144 58106 279290
rect 58274 279144 60314 279290
rect 60482 279144 62522 279290
rect 62690 279144 64730 279290
rect 64898 279144 66938 279290
rect 67106 279144 69146 279290
rect 69314 279144 71354 279290
rect 71522 279144 73562 279290
rect 73730 279144 75770 279290
rect 75938 279144 77978 279290
rect 78146 279144 80186 279290
rect 80354 279144 82394 279290
rect 82562 279144 84602 279290
rect 84770 279144 86810 279290
rect 86978 279144 89018 279290
rect 89186 279144 91226 279290
rect 91394 279144 93434 279290
rect 93602 279144 95642 279290
rect 95810 279144 97850 279290
rect 98018 279144 100058 279290
rect 100226 279144 102266 279290
rect 102434 279144 104474 279290
rect 104642 279144 106682 279290
rect 106850 279144 108890 279290
rect 109058 279144 111098 279290
rect 111266 279144 113306 279290
rect 113474 279144 115514 279290
rect 115682 279144 117722 279290
rect 117890 279144 119930 279290
rect 120098 279144 122138 279290
rect 122306 279144 124346 279290
rect 124514 279144 126554 279290
rect 126722 279144 128762 279290
rect 128930 279144 130970 279290
rect 131138 279144 133178 279290
rect 133346 279144 135386 279290
rect 135554 279144 137594 279290
rect 137762 279144 139802 279290
rect 139970 279144 142010 279290
rect 142178 279144 144218 279290
rect 144386 279144 146426 279290
rect 146594 279144 148634 279290
rect 148802 279144 150842 279290
rect 151010 279144 153050 279290
rect 153218 279144 155258 279290
rect 155426 279144 157466 279290
rect 157634 279144 159674 279290
rect 159842 279144 161882 279290
rect 162050 279144 164090 279290
rect 164258 279144 166298 279290
rect 166466 279144 168506 279290
rect 168674 279144 170714 279290
rect 170882 279144 172922 279290
rect 173090 279144 175130 279290
rect 175298 279144 177338 279290
rect 177506 279144 179546 279290
rect 179714 279144 181754 279290
rect 181922 279144 183962 279290
rect 184130 279144 186170 279290
rect 186338 279144 188378 279290
rect 188546 279144 190586 279290
rect 190754 279144 192794 279290
rect 192962 279144 195002 279290
rect 195170 279144 197210 279290
rect 197378 279144 199418 279290
rect 199586 279144 201626 279290
rect 201794 279144 203834 279290
rect 204002 279144 206042 279290
rect 206210 279144 208250 279290
rect 208418 279144 210458 279290
rect 210626 279144 212666 279290
rect 212834 279144 214874 279290
rect 215042 279144 217082 279290
rect 217250 279144 219290 279290
rect 219458 279144 221498 279290
rect 221666 279144 223706 279290
rect 223874 279144 225914 279290
rect 226082 279144 228122 279290
rect 228290 279144 230330 279290
rect 230498 279144 232538 279290
rect 232706 279144 234746 279290
rect 234914 279144 236954 279290
rect 237122 279144 239162 279290
rect 239330 279144 241370 279290
rect 241538 279144 243578 279290
rect 243746 279144 245786 279290
rect 245954 279144 247994 279290
rect 248162 279144 250202 279290
rect 250370 279144 252410 279290
rect 252578 279144 254618 279290
rect 1676 856 254728 279144
rect 1676 734 16706 856
rect 16874 734 17166 856
rect 17334 734 17626 856
rect 17794 734 18086 856
rect 18254 734 18546 856
rect 18714 734 19006 856
rect 19174 734 19466 856
rect 19634 734 19926 856
rect 20094 734 20386 856
rect 20554 734 20846 856
rect 21014 734 21306 856
rect 21474 734 21766 856
rect 21934 734 22226 856
rect 22394 734 22686 856
rect 22854 734 23146 856
rect 23314 734 23606 856
rect 23774 734 24066 856
rect 24234 734 24526 856
rect 24694 734 24986 856
rect 25154 734 25446 856
rect 25614 734 25906 856
rect 26074 734 26366 856
rect 26534 734 26826 856
rect 26994 734 27286 856
rect 27454 734 27746 856
rect 27914 734 28206 856
rect 28374 734 28666 856
rect 28834 734 29126 856
rect 29294 734 29586 856
rect 29754 734 30046 856
rect 30214 734 30506 856
rect 30674 734 30966 856
rect 31134 734 31426 856
rect 31594 734 31886 856
rect 32054 734 32346 856
rect 32514 734 32806 856
rect 32974 734 33266 856
rect 33434 734 33726 856
rect 33894 734 34186 856
rect 34354 734 34646 856
rect 34814 734 35106 856
rect 35274 734 35566 856
rect 35734 734 36026 856
rect 36194 734 36486 856
rect 36654 734 36946 856
rect 37114 734 37406 856
rect 37574 734 37866 856
rect 38034 734 38326 856
rect 38494 734 38786 856
rect 38954 734 39246 856
rect 39414 734 39706 856
rect 39874 734 40166 856
rect 40334 734 40626 856
rect 40794 734 41086 856
rect 41254 734 41546 856
rect 41714 734 42006 856
rect 42174 734 42466 856
rect 42634 734 42926 856
rect 43094 734 43386 856
rect 43554 734 43846 856
rect 44014 734 44306 856
rect 44474 734 44766 856
rect 44934 734 45226 856
rect 45394 734 45686 856
rect 45854 734 46146 856
rect 46314 734 46606 856
rect 46774 734 47066 856
rect 47234 734 47526 856
rect 47694 734 47986 856
rect 48154 734 48446 856
rect 48614 734 48906 856
rect 49074 734 49366 856
rect 49534 734 49826 856
rect 49994 734 50286 856
rect 50454 734 50746 856
rect 50914 734 51206 856
rect 51374 734 51666 856
rect 51834 734 52126 856
rect 52294 734 52586 856
rect 52754 734 53046 856
rect 53214 734 53506 856
rect 53674 734 53966 856
rect 54134 734 54426 856
rect 54594 734 54886 856
rect 55054 734 55346 856
rect 55514 734 55806 856
rect 55974 734 56266 856
rect 56434 734 56726 856
rect 56894 734 57186 856
rect 57354 734 57646 856
rect 57814 734 58106 856
rect 58274 734 58566 856
rect 58734 734 59026 856
rect 59194 734 59486 856
rect 59654 734 59946 856
rect 60114 734 60406 856
rect 60574 734 60866 856
rect 61034 734 61326 856
rect 61494 734 61786 856
rect 61954 734 62246 856
rect 62414 734 62706 856
rect 62874 734 63166 856
rect 63334 734 63626 856
rect 63794 734 64086 856
rect 64254 734 64546 856
rect 64714 734 65006 856
rect 65174 734 65466 856
rect 65634 734 65926 856
rect 66094 734 66386 856
rect 66554 734 66846 856
rect 67014 734 67306 856
rect 67474 734 67766 856
rect 67934 734 68226 856
rect 68394 734 68686 856
rect 68854 734 69146 856
rect 69314 734 69606 856
rect 69774 734 70066 856
rect 70234 734 70526 856
rect 70694 734 70986 856
rect 71154 734 71446 856
rect 71614 734 71906 856
rect 72074 734 72366 856
rect 72534 734 72826 856
rect 72994 734 73286 856
rect 73454 734 73746 856
rect 73914 734 74206 856
rect 74374 734 74666 856
rect 74834 734 75126 856
rect 75294 734 75586 856
rect 75754 734 76046 856
rect 76214 734 76506 856
rect 76674 734 76966 856
rect 77134 734 77426 856
rect 77594 734 77886 856
rect 78054 734 78346 856
rect 78514 734 78806 856
rect 78974 734 79266 856
rect 79434 734 79726 856
rect 79894 734 80186 856
rect 80354 734 80646 856
rect 80814 734 81106 856
rect 81274 734 81566 856
rect 81734 734 82026 856
rect 82194 734 82486 856
rect 82654 734 82946 856
rect 83114 734 83406 856
rect 83574 734 83866 856
rect 84034 734 84326 856
rect 84494 734 84786 856
rect 84954 734 85246 856
rect 85414 734 85706 856
rect 85874 734 86166 856
rect 86334 734 86626 856
rect 86794 734 87086 856
rect 87254 734 87546 856
rect 87714 734 88006 856
rect 88174 734 88466 856
rect 88634 734 88926 856
rect 89094 734 89386 856
rect 89554 734 89846 856
rect 90014 734 90306 856
rect 90474 734 90766 856
rect 90934 734 91226 856
rect 91394 734 91686 856
rect 91854 734 92146 856
rect 92314 734 92606 856
rect 92774 734 93066 856
rect 93234 734 93526 856
rect 93694 734 93986 856
rect 94154 734 94446 856
rect 94614 734 94906 856
rect 95074 734 95366 856
rect 95534 734 95826 856
rect 95994 734 96286 856
rect 96454 734 96746 856
rect 96914 734 97206 856
rect 97374 734 97666 856
rect 97834 734 98126 856
rect 98294 734 98586 856
rect 98754 734 99046 856
rect 99214 734 99506 856
rect 99674 734 99966 856
rect 100134 734 100426 856
rect 100594 734 100886 856
rect 101054 734 101346 856
rect 101514 734 101806 856
rect 101974 734 102266 856
rect 102434 734 102726 856
rect 102894 734 103186 856
rect 103354 734 103646 856
rect 103814 734 104106 856
rect 104274 734 104566 856
rect 104734 734 105026 856
rect 105194 734 105486 856
rect 105654 734 105946 856
rect 106114 734 106406 856
rect 106574 734 106866 856
rect 107034 734 107326 856
rect 107494 734 107786 856
rect 107954 734 108246 856
rect 108414 734 108706 856
rect 108874 734 109166 856
rect 109334 734 109626 856
rect 109794 734 110086 856
rect 110254 734 110546 856
rect 110714 734 111006 856
rect 111174 734 111466 856
rect 111634 734 111926 856
rect 112094 734 112386 856
rect 112554 734 112846 856
rect 113014 734 113306 856
rect 113474 734 113766 856
rect 113934 734 114226 856
rect 114394 734 114686 856
rect 114854 734 115146 856
rect 115314 734 115606 856
rect 115774 734 116066 856
rect 116234 734 116526 856
rect 116694 734 116986 856
rect 117154 734 117446 856
rect 117614 734 117906 856
rect 118074 734 118366 856
rect 118534 734 118826 856
rect 118994 734 119286 856
rect 119454 734 119746 856
rect 119914 734 120206 856
rect 120374 734 120666 856
rect 120834 734 121126 856
rect 121294 734 121586 856
rect 121754 734 122046 856
rect 122214 734 122506 856
rect 122674 734 122966 856
rect 123134 734 123426 856
rect 123594 734 123886 856
rect 124054 734 124346 856
rect 124514 734 124806 856
rect 124974 734 125266 856
rect 125434 734 125726 856
rect 125894 734 126186 856
rect 126354 734 126646 856
rect 126814 734 127106 856
rect 127274 734 127566 856
rect 127734 734 128026 856
rect 128194 734 128486 856
rect 128654 734 128946 856
rect 129114 734 129406 856
rect 129574 734 129866 856
rect 130034 734 130326 856
rect 130494 734 130786 856
rect 130954 734 131246 856
rect 131414 734 131706 856
rect 131874 734 132166 856
rect 132334 734 132626 856
rect 132794 734 133086 856
rect 133254 734 133546 856
rect 133714 734 134006 856
rect 134174 734 134466 856
rect 134634 734 134926 856
rect 135094 734 135386 856
rect 135554 734 135846 856
rect 136014 734 136306 856
rect 136474 734 136766 856
rect 136934 734 137226 856
rect 137394 734 137686 856
rect 137854 734 138146 856
rect 138314 734 138606 856
rect 138774 734 139066 856
rect 139234 734 139526 856
rect 139694 734 139986 856
rect 140154 734 140446 856
rect 140614 734 140906 856
rect 141074 734 141366 856
rect 141534 734 141826 856
rect 141994 734 142286 856
rect 142454 734 142746 856
rect 142914 734 143206 856
rect 143374 734 143666 856
rect 143834 734 144126 856
rect 144294 734 144586 856
rect 144754 734 145046 856
rect 145214 734 145506 856
rect 145674 734 145966 856
rect 146134 734 146426 856
rect 146594 734 146886 856
rect 147054 734 147346 856
rect 147514 734 147806 856
rect 147974 734 148266 856
rect 148434 734 148726 856
rect 148894 734 149186 856
rect 149354 734 149646 856
rect 149814 734 150106 856
rect 150274 734 150566 856
rect 150734 734 151026 856
rect 151194 734 151486 856
rect 151654 734 151946 856
rect 152114 734 152406 856
rect 152574 734 152866 856
rect 153034 734 153326 856
rect 153494 734 153786 856
rect 153954 734 154246 856
rect 154414 734 154706 856
rect 154874 734 155166 856
rect 155334 734 155626 856
rect 155794 734 156086 856
rect 156254 734 156546 856
rect 156714 734 157006 856
rect 157174 734 157466 856
rect 157634 734 157926 856
rect 158094 734 158386 856
rect 158554 734 158846 856
rect 159014 734 159306 856
rect 159474 734 159766 856
rect 159934 734 160226 856
rect 160394 734 160686 856
rect 160854 734 161146 856
rect 161314 734 161606 856
rect 161774 734 162066 856
rect 162234 734 162526 856
rect 162694 734 162986 856
rect 163154 734 163446 856
rect 163614 734 163906 856
rect 164074 734 164366 856
rect 164534 734 164826 856
rect 164994 734 165286 856
rect 165454 734 165746 856
rect 165914 734 166206 856
rect 166374 734 166666 856
rect 166834 734 167126 856
rect 167294 734 167586 856
rect 167754 734 168046 856
rect 168214 734 168506 856
rect 168674 734 168966 856
rect 169134 734 169426 856
rect 169594 734 169886 856
rect 170054 734 170346 856
rect 170514 734 170806 856
rect 170974 734 171266 856
rect 171434 734 171726 856
rect 171894 734 172186 856
rect 172354 734 172646 856
rect 172814 734 173106 856
rect 173274 734 173566 856
rect 173734 734 174026 856
rect 174194 734 174486 856
rect 174654 734 174946 856
rect 175114 734 175406 856
rect 175574 734 175866 856
rect 176034 734 176326 856
rect 176494 734 176786 856
rect 176954 734 177246 856
rect 177414 734 177706 856
rect 177874 734 178166 856
rect 178334 734 178626 856
rect 178794 734 179086 856
rect 179254 734 179546 856
rect 179714 734 180006 856
rect 180174 734 180466 856
rect 180634 734 180926 856
rect 181094 734 181386 856
rect 181554 734 181846 856
rect 182014 734 182306 856
rect 182474 734 182766 856
rect 182934 734 183226 856
rect 183394 734 183686 856
rect 183854 734 184146 856
rect 184314 734 184606 856
rect 184774 734 185066 856
rect 185234 734 185526 856
rect 185694 734 185986 856
rect 186154 734 186446 856
rect 186614 734 186906 856
rect 187074 734 187366 856
rect 187534 734 187826 856
rect 187994 734 188286 856
rect 188454 734 188746 856
rect 188914 734 189206 856
rect 189374 734 189666 856
rect 189834 734 190126 856
rect 190294 734 190586 856
rect 190754 734 191046 856
rect 191214 734 191506 856
rect 191674 734 191966 856
rect 192134 734 192426 856
rect 192594 734 192886 856
rect 193054 734 193346 856
rect 193514 734 193806 856
rect 193974 734 194266 856
rect 194434 734 194726 856
rect 194894 734 195186 856
rect 195354 734 195646 856
rect 195814 734 196106 856
rect 196274 734 196566 856
rect 196734 734 197026 856
rect 197194 734 197486 856
rect 197654 734 197946 856
rect 198114 734 198406 856
rect 198574 734 198866 856
rect 199034 734 199326 856
rect 199494 734 199786 856
rect 199954 734 200246 856
rect 200414 734 200706 856
rect 200874 734 201166 856
rect 201334 734 201626 856
rect 201794 734 202086 856
rect 202254 734 202546 856
rect 202714 734 203006 856
rect 203174 734 203466 856
rect 203634 734 203926 856
rect 204094 734 204386 856
rect 204554 734 204846 856
rect 205014 734 205306 856
rect 205474 734 205766 856
rect 205934 734 206226 856
rect 206394 734 206686 856
rect 206854 734 207146 856
rect 207314 734 207606 856
rect 207774 734 208066 856
rect 208234 734 208526 856
rect 208694 734 208986 856
rect 209154 734 209446 856
rect 209614 734 209906 856
rect 210074 734 210366 856
rect 210534 734 210826 856
rect 210994 734 211286 856
rect 211454 734 211746 856
rect 211914 734 212206 856
rect 212374 734 212666 856
rect 212834 734 213126 856
rect 213294 734 213586 856
rect 213754 734 214046 856
rect 214214 734 214506 856
rect 214674 734 214966 856
rect 215134 734 215426 856
rect 215594 734 215886 856
rect 216054 734 216346 856
rect 216514 734 216806 856
rect 216974 734 217266 856
rect 217434 734 217726 856
rect 217894 734 218186 856
rect 218354 734 218646 856
rect 218814 734 219106 856
rect 219274 734 219566 856
rect 219734 734 220026 856
rect 220194 734 220486 856
rect 220654 734 220946 856
rect 221114 734 221406 856
rect 221574 734 221866 856
rect 222034 734 222326 856
rect 222494 734 222786 856
rect 222954 734 223246 856
rect 223414 734 223706 856
rect 223874 734 224166 856
rect 224334 734 224626 856
rect 224794 734 225086 856
rect 225254 734 225546 856
rect 225714 734 226006 856
rect 226174 734 226466 856
rect 226634 734 226926 856
rect 227094 734 227386 856
rect 227554 734 227846 856
rect 228014 734 228306 856
rect 228474 734 228766 856
rect 228934 734 229226 856
rect 229394 734 229686 856
rect 229854 734 230146 856
rect 230314 734 230606 856
rect 230774 734 231066 856
rect 231234 734 231526 856
rect 231694 734 231986 856
rect 232154 734 232446 856
rect 232614 734 232906 856
rect 233074 734 233366 856
rect 233534 734 233826 856
rect 233994 734 234286 856
rect 234454 734 234746 856
rect 234914 734 235206 856
rect 235374 734 235666 856
rect 235834 734 236126 856
rect 236294 734 236586 856
rect 236754 734 237046 856
rect 237214 734 237506 856
rect 237674 734 237966 856
rect 238134 734 238426 856
rect 238594 734 238886 856
rect 239054 734 239346 856
rect 239514 734 239806 856
rect 239974 734 240266 856
rect 240434 734 240726 856
rect 240894 734 241186 856
rect 241354 734 241646 856
rect 241814 734 242106 856
rect 242274 734 242566 856
rect 242734 734 243026 856
rect 243194 734 254728 856
<< obsm3 >>
rect 2313 2143 250286 277473
<< metal4 >>
rect 4208 2128 4528 277488
rect 19568 2128 19888 277488
rect 34928 2128 35248 277488
rect 50288 2128 50608 277488
rect 65648 2128 65968 277488
rect 81008 2128 81328 277488
rect 96368 2128 96688 277488
rect 111728 2128 112048 277488
rect 127088 2128 127408 277488
rect 142448 2128 142768 277488
rect 157808 2128 158128 277488
rect 173168 2128 173488 277488
rect 188528 2128 188848 277488
rect 203888 2128 204208 277488
rect 219248 2128 219568 277488
rect 234608 2128 234928 277488
rect 249968 2128 250288 277488
<< obsm4 >>
rect 3187 2211 4128 277133
rect 4608 2211 19488 277133
rect 19968 2211 34848 277133
rect 35328 2211 50208 277133
rect 50688 2211 65568 277133
rect 66048 2211 80928 277133
rect 81408 2211 96288 277133
rect 96768 2211 111648 277133
rect 112128 2211 127008 277133
rect 127488 2211 142368 277133
rect 142848 2211 157728 277133
rect 158208 2211 173088 277133
rect 173568 2211 188448 277133
rect 188928 2211 203808 277133
rect 204288 2211 219168 277133
rect 219648 2211 223869 277133
<< labels >>
rlabel metal2 s 5170 279200 5226 280000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 71410 279200 71466 280000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 78034 279200 78090 280000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 84658 279200 84714 280000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 91282 279200 91338 280000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 97906 279200 97962 280000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 104530 279200 104586 280000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 111154 279200 111210 280000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 117778 279200 117834 280000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 124402 279200 124458 280000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 131026 279200 131082 280000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 11794 279200 11850 280000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 137650 279200 137706 280000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 144274 279200 144330 280000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 150898 279200 150954 280000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 157522 279200 157578 280000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 164146 279200 164202 280000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 170770 279200 170826 280000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 177394 279200 177450 280000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 184018 279200 184074 280000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 190642 279200 190698 280000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 197266 279200 197322 280000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 18418 279200 18474 280000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 203890 279200 203946 280000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 210514 279200 210570 280000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 217138 279200 217194 280000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 223762 279200 223818 280000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 230386 279200 230442 280000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 237010 279200 237066 280000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 243634 279200 243690 280000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 250258 279200 250314 280000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 25042 279200 25098 280000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 31666 279200 31722 280000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 38290 279200 38346 280000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 44914 279200 44970 280000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 51538 279200 51594 280000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 58162 279200 58218 280000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 64786 279200 64842 280000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 7378 279200 7434 280000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 73618 279200 73674 280000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 80242 279200 80298 280000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 86866 279200 86922 280000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 93490 279200 93546 280000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 100114 279200 100170 280000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 106738 279200 106794 280000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 113362 279200 113418 280000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 119986 279200 120042 280000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 126610 279200 126666 280000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 133234 279200 133290 280000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 14002 279200 14058 280000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 139858 279200 139914 280000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 146482 279200 146538 280000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 153106 279200 153162 280000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 159730 279200 159786 280000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 166354 279200 166410 280000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 172978 279200 173034 280000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 179602 279200 179658 280000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 186226 279200 186282 280000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 192850 279200 192906 280000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 199474 279200 199530 280000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 20626 279200 20682 280000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 206098 279200 206154 280000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 212722 279200 212778 280000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 219346 279200 219402 280000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 225970 279200 226026 280000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 232594 279200 232650 280000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 239218 279200 239274 280000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 245842 279200 245898 280000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 252466 279200 252522 280000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 27250 279200 27306 280000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 33874 279200 33930 280000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 40498 279200 40554 280000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 47122 279200 47178 280000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 53746 279200 53802 280000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 60370 279200 60426 280000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 66994 279200 67050 280000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9586 279200 9642 280000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 75826 279200 75882 280000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 82450 279200 82506 280000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 89074 279200 89130 280000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 95698 279200 95754 280000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 102322 279200 102378 280000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 108946 279200 109002 280000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 115570 279200 115626 280000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 122194 279200 122250 280000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 128818 279200 128874 280000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 135442 279200 135498 280000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 16210 279200 16266 280000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 142066 279200 142122 280000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 148690 279200 148746 280000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 155314 279200 155370 280000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 161938 279200 161994 280000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 168562 279200 168618 280000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 175186 279200 175242 280000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 181810 279200 181866 280000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 188434 279200 188490 280000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 195058 279200 195114 280000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 201682 279200 201738 280000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 22834 279200 22890 280000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 208306 279200 208362 280000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 214930 279200 214986 280000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 221554 279200 221610 280000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 228178 279200 228234 280000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 234802 279200 234858 280000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 241426 279200 241482 280000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 248050 279200 248106 280000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 254674 279200 254730 280000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 29458 279200 29514 280000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 36082 279200 36138 280000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 42706 279200 42762 280000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 49330 279200 49386 280000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 55954 279200 56010 280000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 62578 279200 62634 280000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 69202 279200 69258 280000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 242162 0 242218 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 242622 0 242678 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 243082 0 243138 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 203522 0 203578 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 204902 0 204958 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 209042 0 209098 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 221462 0 221518 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 224222 0 224278 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 225602 0 225658 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 226982 0 227038 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 231122 0 231178 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 238022 0 238078 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 151082 0 151138 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 163502 0 163558 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 170402 0 170458 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 180062 0 180118 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 181442 0 181498 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 189722 0 189778 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 196622 0 196678 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 205362 0 205418 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 208122 0 208178 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 209502 0 209558 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 212262 0 212318 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 213642 0 213698 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 217782 0 217838 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 220542 0 220598 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 221922 0 221978 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 223302 0 223358 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 224682 0 224738 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 226062 0 226118 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 227442 0 227498 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 228822 0 228878 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 230202 0 230258 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 231582 0 231638 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 232962 0 233018 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 234342 0 234398 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 235722 0 235778 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 237102 0 237158 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 238482 0 238538 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 239862 0 239918 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 241242 0 241298 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 121182 0 121238 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 144642 0 144698 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 147402 0 147458 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 155682 0 155738 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 159822 0 159878 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 165342 0 165398 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 168102 0 168158 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 177762 0 177818 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 180522 0 180578 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 183282 0 183338 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 186042 0 186098 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 190182 0 190238 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 191562 0 191618 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 192942 0 192998 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 195702 0 195758 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 198462 0 198518 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 199842 0 199898 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 201222 0 201278 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 202602 0 202658 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 204442 0 204498 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 212722 0 212778 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 214102 0 214158 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 215482 0 215538 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 216862 0 216918 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 219622 0 219678 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 223762 0 223818 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 227902 0 227958 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 236182 0 236238 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 240322 0 240378 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 241702 0 241758 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 182362 0 182418 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 189262 0 189318 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 200302 0 200358 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 201682 0 201738 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 277488 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 277488 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 16762 0 16818 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 260000 280000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 146014906
string GDS_FILE /si/work/caravel-gf180-pio/openlane/wb_pio/runs/sky130B-2022-12-28_12_25/results/signoff/wb_pio.magic.gds
string GDS_START 1332350
<< end >>

